//Copyright (C)2014-2024 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: Post-PnR Verilog Simulation Model file
//Tool Version: V1.9.10.03 Education
//Created Time: Sat May 10 14:52:18 2025

`timescale 100 ps/100 ps
module SDRAM_Controller_HS_Top(
	I_sdrc_rst_n,
	I_sdrc_clk,
	I_sdram_clk,
	I_sdrc_cmd_en,
	I_sdrc_cmd,
	I_sdrc_precharge_ctrl,
	I_sdram_power_down,
	I_sdram_selfrefresh,
	I_sdrc_addr,
	I_sdrc_dqm,
	I_sdrc_data,
	I_sdrc_data_len,
	O_sdram_clk,
	O_sdram_cke,
	O_sdram_cs_n,
	O_sdram_cas_n,
	O_sdram_ras_n,
	O_sdram_wen_n,
	O_sdram_dqm,
	O_sdram_addr,
	O_sdram_ba,
	O_sdrc_data,
	O_sdrc_init_done,
	O_sdrc_cmd_ack,
	IO_sdram_dq
);
input I_sdrc_rst_n;
input I_sdrc_clk;
input I_sdram_clk;
input I_sdrc_cmd_en;
input [2:0] I_sdrc_cmd;
input I_sdrc_precharge_ctrl;
input I_sdram_power_down;
input I_sdram_selfrefresh;
input [20:0] I_sdrc_addr;
input [3:0] I_sdrc_dqm;
input [31:0] I_sdrc_data;
input [7:0] I_sdrc_data_len;
output O_sdram_clk;
output O_sdram_cke;
output O_sdram_cs_n;
output O_sdram_cas_n;
output O_sdram_ras_n;
output O_sdram_wen_n;
output [3:0] O_sdram_dqm;
output [10:0] O_sdram_addr;
output [1:0] O_sdram_ba;
output [31:0] O_sdrc_data;
output O_sdrc_init_done;
output O_sdrc_cmd_ack;
inout [31:0] IO_sdram_dq;
wire [31:0] Ctrl_fsm_data;
wire GND;
wire [31:0] IO_sdram_dq;
wire IO_sdram_dq_0_6;
wire [31:0] IO_sdram_dq_in;
wire I_sdram_clk;
wire I_sdram_power_down;
wire I_sdram_selfrefresh;
wire [20:0] I_sdrc_addr;
wire I_sdrc_clk;
wire [2:0] I_sdrc_cmd;
wire I_sdrc_cmd_en;
wire [31:0] I_sdrc_data;
wire [7:0] I_sdrc_data_len;
wire [3:0] I_sdrc_dqm;
wire I_sdrc_precharge_ctrl;
wire I_sdrc_rst_n;
wire [10:0] O_sdram_addr;
wire [1:0] O_sdram_ba;
wire O_sdram_cas_n;
wire O_sdram_cke;
wire O_sdram_clk;
wire O_sdram_cs_n;
wire [3:0] O_sdram_dqm;
wire O_sdram_ras_n;
wire O_sdram_wen_n;
wire O_sdrc_cmd_ack;
wire [31:0] O_sdrc_data;
wire O_sdrc_init_done;
wire VCC;
wire \u_sdrc_hs_top/n202_5 ;
wire \u_sdrc_hs_top/n204_5 ;
wire \u_sdrc_hs_top/n153_15 ;
wire \u_sdrc_hs_top/n155_16 ;
wire \u_sdrc_hs_top/n157_16 ;
wire \u_sdrc_hs_top/n159_16 ;
wire \u_sdrc_hs_top/n161_15 ;
wire \u_sdrc_hs_top/n163_16 ;
wire \u_sdrc_hs_top/n169_16 ;
wire \u_sdrc_hs_top/n171_17 ;
wire \u_sdrc_hs_top/n65_4 ;
wire \u_sdrc_hs_top/n64_4 ;
wire \u_sdrc_hs_top/n63_4 ;
wire \u_sdrc_hs_top/n153_16 ;
wire \u_sdrc_hs_top/n155_17 ;
wire \u_sdrc_hs_top/n157_17 ;
wire \u_sdrc_hs_top/n163_17 ;
wire \u_sdrc_hs_top/n153_17 ;
wire \u_sdrc_hs_top/n163_18 ;
wire \u_sdrc_hs_top/n167_18 ;
wire \u_sdrc_hs_top/n165_19 ;
wire \u_sdrc_hs_top/n200_7 ;
wire \u_sdrc_hs_top/n27_11 ;
wire \u_sdrc_hs_top/n67_6 ;
wire \u_sdrc_hs_top/Cmd_init_state.INIT_STATE_PRECHARGEALL ;
wire \u_sdrc_hs_top/Cmd_init_state.INIT_STATE_AUTOREFRESH1 ;
wire \u_sdrc_hs_top/Cmd_init_state.INIT_STATE_AUTOREFRESH2 ;
wire \u_sdrc_hs_top/Cmd_init_state.INIT_STATE_LOAD_MODEREG ;
wire \u_sdrc_hs_top/Cmd_init_state.INIT_STATE_PRECHARGE_DELAY ;
wire \u_sdrc_hs_top/Cmd_init_state.INIT_STATE_AUTOREFRESH1_DELAY ;
wire \u_sdrc_hs_top/Cmd_init_state.INIT_STATE_AUTOREFRESH2_DELAY ;
wire \u_sdrc_hs_top/Cmd_init_state.INIT_STATE_LOAD_MODEREG_DELAY ;
wire \u_sdrc_hs_top/Cmd_init_state.INIT_STATE_INIT_DONE ;
wire \u_sdrc_hs_top/Cmd_init_state.INIT_STATE_IDLE ;
wire \u_sdrc_hs_top/U_ODDR_clk_1_Q1 ;
wire \u_sdrc_hs_top/n26_1 ;
wire \u_sdrc_hs_top/n26_2 ;
wire \u_sdrc_hs_top/n25_1 ;
wire \u_sdrc_hs_top/n25_2 ;
wire \u_sdrc_hs_top/n24_1 ;
wire \u_sdrc_hs_top/n24_2 ;
wire \u_sdrc_hs_top/n23_1 ;
wire \u_sdrc_hs_top/n23_2 ;
wire \u_sdrc_hs_top/n22_1 ;
wire \u_sdrc_hs_top/n22_2 ;
wire \u_sdrc_hs_top/n21_1 ;
wire \u_sdrc_hs_top/n21_2 ;
wire \u_sdrc_hs_top/n20_1 ;
wire \u_sdrc_hs_top/n20_2 ;
wire \u_sdrc_hs_top/n19_1 ;
wire \u_sdrc_hs_top/n19_2 ;
wire \u_sdrc_hs_top/n18_1 ;
wire \u_sdrc_hs_top/n18_2 ;
wire \u_sdrc_hs_top/n17_1 ;
wire \u_sdrc_hs_top/n17_2 ;
wire \u_sdrc_hs_top/n16_1 ;
wire \u_sdrc_hs_top/n16_2 ;
wire \u_sdrc_hs_top/n15_1 ;
wire \u_sdrc_hs_top/n15_2 ;
wire \u_sdrc_hs_top/n14_1 ;
wire \u_sdrc_hs_top/n14_2 ;
wire \u_sdrc_hs_top/n13_1 ;
wire \u_sdrc_hs_top/n13_2 ;
wire \u_sdrc_hs_top/n12_1 ;
wire \u_sdrc_hs_top/n12_0_COUT ;
wire \u_sdrc_hs_top/n9_6 ;
wire \u_sdrc_hs_top/n205_6 ;
wire \u_sdrc_hs_top/n66_6 ;
wire \u_sdrc_hs_top/Init_cnt_14_9 ;
wire \u_sdrc_hs_top/Sdram_wen_n ;
wire \u_sdrc_hs_top/Sdram_cas_n ;
wire \u_sdrc_hs_top/Sdram_ras_n ;
wire \u_sdrc_hs_top/Sdram_cke ;
wire [15:0] \u_sdrc_hs_top/Init_cnt ;
wire [3:0] \u_sdrc_hs_top/Count_init_delay ;
wire [2:0] \u_sdrc_hs_top/Sdram_cmd_init ;
wire [1:1] \u_sdrc_hs_top/Sdram_ba_init ;
wire [1:0] \u_sdrc_hs_top/Sdram_ba ;
wire [10:0] \u_sdrc_hs_top/Sdram_addr ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n179_3 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n180_3 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n181_3 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n182_3 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n183_3 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n184_3 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n185_3 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n186_3 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_wr_data_valid_8 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n80_29 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n590_31 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n592_31 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n997_16 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1003_16 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n580_32 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n582_31 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n584_32 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n586_31 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n588_31 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n594_31 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n596_33 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n598_33 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n602_32 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n604_31 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1000_17 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1005_18 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1007_18 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1009_18 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1011_18 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1013_18 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1015_18 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1017_18 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1019_18 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1021_18 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1023_18 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1025_18 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1027_18 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1029_18 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n80_31 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n606_14 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n618_12 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_cke_7 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n86_4 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n85_4 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n84_4 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n100_4 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n99_4 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n98_4 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n179_4 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n179_5 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n181_5 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n182_4 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n182_5 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n183_5 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n184_4 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n184_5 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n185_4 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n993_4 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd_7_9 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_wr_data_valid_9 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n80_32 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n590_32 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n590_33 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n592_33 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n592_35 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n997_17 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n997_18 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1003_17 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1003_18 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n582_32 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n582_33 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n582_34 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n582_35 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n584_33 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n586_32 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n586_33 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n588_32 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n598_34 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1000_18 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1000_19 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1005_19 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1005_20 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1005_21 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1007_19 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1007_20 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1009_20 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1011_19 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1013_19 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1015_19 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1015_20 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1017_19 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1017_20 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1019_19 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1019_20 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1021_19 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1021_20 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1023_19 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1023_20 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1025_19 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1025_20 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1027_19 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1027_20 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1029_19 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1029_20 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n80_33 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n80_34 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n614_13 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n616_13 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n759_6 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_cke_8 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n181_6 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n993_5 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_wr_data_valid_10 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_wr_data_valid_11 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_wr_data_valid_12 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n590_34 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n592_36 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n997_19 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n997_20 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1003_19 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1003_20 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1003_22 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n582_36 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n582_38 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n582_39 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n582_40 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n582_41 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n582_42 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n586_34 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n598_35 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1000_20 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1000_21 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1005_22 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1007_21 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1007_22 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1009_21 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1011_20 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1013_20 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1015_21 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1017_21 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1019_21 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1021_21 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1023_21 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1025_21 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1027_21 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1029_21 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n80_35 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_wr_data_valid_13 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_wr_data_valid_14 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n590_35 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1003_23 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n582_43 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n582_44 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n582_45 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n582_46 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n582_47 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n582_49 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n582_50 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1000_22 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1005_23 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1005_24 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1009_22 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1015_22 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1017_22 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1019_22 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1019_23 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1021_22 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1023_22 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1025_22 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1027_22 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1029_22 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n997_22 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n181_8 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n180_8 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n179_8 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n183_7 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n592_38 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n610_15 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n612_15 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n582_52 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n993_7 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n584_36 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n580_36 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/Reset_cmd_count ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1003_25 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n759_8 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n997_24 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n582_54 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n1009_24 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n80_38 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n592_40 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n620_14 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n616_15 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n614_15 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n610_17 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n608_14 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd_7_11 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n622_17 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n606_17 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n180_10 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n606_19 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n580_38 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/Precharge_flag ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_AUTOREFRESH_DELAY ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_IDLE ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_ACTIVE2RW_DELAY ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_READ_WITHOUT_AUTOPRE ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_WRITE_WITHOUT_AUTOPRE ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_DATAIN2ACTIVE ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_PRECHARGE_DELAY ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_INIT ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_POWER_DOWN ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_SELFREFRESH ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_SELFREFRESH_WAIT ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_SELFREFRESH_EXIT ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_wr_data_valid ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n87_6 ;
wire \u_sdrc_hs_top/u_sdrc_control_fsm/n101_6 ;
wire [3:0] \u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay ;
wire [3:0] \u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay2 ;
wire [7:0] \u_sdrc_hs_top/u_sdrc_control_fsm/Sdrc_wrd_len ;
wire [1:0] \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_bk_wrd ;
wire [7:0] \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd ;
wire [8:0] \u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num ;
VCC VCC_cZ (
  .V(VCC)
);
GND GND_cZ (
  .G(GND)
);
// GSR GSR (
// 	.GSRI(VCC)
// );
IOBUF IO_sdram_dq_0_iobuf (
	.I(Ctrl_fsm_data[0]),
	.OEN(IO_sdram_dq_0_6),
	.IO(IO_sdram_dq[0]),
	.O(IO_sdram_dq_in[0])
);
IOBUF IO_sdram_dq_1_iobuf (
	.I(Ctrl_fsm_data[1]),
	.OEN(IO_sdram_dq_0_6),
	.IO(IO_sdram_dq[1]),
	.O(IO_sdram_dq_in[1])
);
IOBUF IO_sdram_dq_2_iobuf (
	.I(Ctrl_fsm_data[2]),
	.OEN(IO_sdram_dq_0_6),
	.IO(IO_sdram_dq[2]),
	.O(IO_sdram_dq_in[2])
);
IOBUF IO_sdram_dq_3_iobuf (
	.I(Ctrl_fsm_data[3]),
	.OEN(IO_sdram_dq_0_6),
	.IO(IO_sdram_dq[3]),
	.O(IO_sdram_dq_in[3])
);
IOBUF IO_sdram_dq_4_iobuf (
	.I(Ctrl_fsm_data[4]),
	.OEN(IO_sdram_dq_0_6),
	.IO(IO_sdram_dq[4]),
	.O(IO_sdram_dq_in[4])
);
IOBUF IO_sdram_dq_5_iobuf (
	.I(Ctrl_fsm_data[5]),
	.OEN(IO_sdram_dq_0_6),
	.IO(IO_sdram_dq[5]),
	.O(IO_sdram_dq_in[5])
);
IOBUF IO_sdram_dq_6_iobuf (
	.I(Ctrl_fsm_data[6]),
	.OEN(IO_sdram_dq_0_6),
	.IO(IO_sdram_dq[6]),
	.O(IO_sdram_dq_in[6])
);
IOBUF IO_sdram_dq_7_iobuf (
	.I(Ctrl_fsm_data[7]),
	.OEN(IO_sdram_dq_0_6),
	.IO(IO_sdram_dq[7]),
	.O(IO_sdram_dq_in[7])
);
IOBUF IO_sdram_dq_8_iobuf (
	.I(Ctrl_fsm_data[8]),
	.OEN(IO_sdram_dq_0_6),
	.IO(IO_sdram_dq[8]),
	.O(IO_sdram_dq_in[8])
);
IOBUF IO_sdram_dq_9_iobuf (
	.I(Ctrl_fsm_data[9]),
	.OEN(IO_sdram_dq_0_6),
	.IO(IO_sdram_dq[9]),
	.O(IO_sdram_dq_in[9])
);
IOBUF IO_sdram_dq_10_iobuf (
	.I(Ctrl_fsm_data[10]),
	.OEN(IO_sdram_dq_0_6),
	.IO(IO_sdram_dq[10]),
	.O(IO_sdram_dq_in[10])
);
IOBUF IO_sdram_dq_11_iobuf (
	.I(Ctrl_fsm_data[11]),
	.OEN(IO_sdram_dq_0_6),
	.IO(IO_sdram_dq[11]),
	.O(IO_sdram_dq_in[11])
);
IOBUF IO_sdram_dq_12_iobuf (
	.I(Ctrl_fsm_data[12]),
	.OEN(IO_sdram_dq_0_6),
	.IO(IO_sdram_dq[12]),
	.O(IO_sdram_dq_in[12])
);
IOBUF IO_sdram_dq_13_iobuf (
	.I(Ctrl_fsm_data[13]),
	.OEN(IO_sdram_dq_0_6),
	.IO(IO_sdram_dq[13]),
	.O(IO_sdram_dq_in[13])
);
IOBUF IO_sdram_dq_14_iobuf (
	.I(Ctrl_fsm_data[14]),
	.OEN(IO_sdram_dq_0_6),
	.IO(IO_sdram_dq[14]),
	.O(IO_sdram_dq_in[14])
);
IOBUF IO_sdram_dq_15_iobuf (
	.I(Ctrl_fsm_data[15]),
	.OEN(IO_sdram_dq_0_6),
	.IO(IO_sdram_dq[15]),
	.O(IO_sdram_dq_in[15])
);
IOBUF IO_sdram_dq_16_iobuf (
	.I(Ctrl_fsm_data[16]),
	.OEN(IO_sdram_dq_0_6),
	.IO(IO_sdram_dq[16]),
	.O(IO_sdram_dq_in[16])
);
IOBUF IO_sdram_dq_17_iobuf (
	.I(Ctrl_fsm_data[17]),
	.OEN(IO_sdram_dq_0_6),
	.IO(IO_sdram_dq[17]),
	.O(IO_sdram_dq_in[17])
);
IOBUF IO_sdram_dq_18_iobuf (
	.I(Ctrl_fsm_data[18]),
	.OEN(IO_sdram_dq_0_6),
	.IO(IO_sdram_dq[18]),
	.O(IO_sdram_dq_in[18])
);
IOBUF IO_sdram_dq_19_iobuf (
	.I(Ctrl_fsm_data[19]),
	.OEN(IO_sdram_dq_0_6),
	.IO(IO_sdram_dq[19]),
	.O(IO_sdram_dq_in[19])
);
IOBUF IO_sdram_dq_20_iobuf (
	.I(Ctrl_fsm_data[20]),
	.OEN(IO_sdram_dq_0_6),
	.IO(IO_sdram_dq[20]),
	.O(IO_sdram_dq_in[20])
);
IOBUF IO_sdram_dq_21_iobuf (
	.I(Ctrl_fsm_data[21]),
	.OEN(IO_sdram_dq_0_6),
	.IO(IO_sdram_dq[21]),
	.O(IO_sdram_dq_in[21])
);
IOBUF IO_sdram_dq_22_iobuf (
	.I(Ctrl_fsm_data[22]),
	.OEN(IO_sdram_dq_0_6),
	.IO(IO_sdram_dq[22]),
	.O(IO_sdram_dq_in[22])
);
IOBUF IO_sdram_dq_23_iobuf (
	.I(Ctrl_fsm_data[23]),
	.OEN(IO_sdram_dq_0_6),
	.IO(IO_sdram_dq[23]),
	.O(IO_sdram_dq_in[23])
);
IOBUF IO_sdram_dq_24_iobuf (
	.I(Ctrl_fsm_data[24]),
	.OEN(IO_sdram_dq_0_6),
	.IO(IO_sdram_dq[24]),
	.O(IO_sdram_dq_in[24])
);
IOBUF IO_sdram_dq_25_iobuf (
	.I(Ctrl_fsm_data[25]),
	.OEN(IO_sdram_dq_0_6),
	.IO(IO_sdram_dq[25]),
	.O(IO_sdram_dq_in[25])
);
IOBUF IO_sdram_dq_26_iobuf (
	.I(Ctrl_fsm_data[26]),
	.OEN(IO_sdram_dq_0_6),
	.IO(IO_sdram_dq[26]),
	.O(IO_sdram_dq_in[26])
);
IOBUF IO_sdram_dq_27_iobuf (
	.I(Ctrl_fsm_data[27]),
	.OEN(IO_sdram_dq_0_6),
	.IO(IO_sdram_dq[27]),
	.O(IO_sdram_dq_in[27])
);
IOBUF IO_sdram_dq_28_iobuf (
	.I(Ctrl_fsm_data[28]),
	.OEN(IO_sdram_dq_0_6),
	.IO(IO_sdram_dq[28]),
	.O(IO_sdram_dq_in[28])
);
IOBUF IO_sdram_dq_29_iobuf (
	.I(Ctrl_fsm_data[29]),
	.OEN(IO_sdram_dq_0_6),
	.IO(IO_sdram_dq[29]),
	.O(IO_sdram_dq_in[29])
);
IOBUF IO_sdram_dq_30_iobuf (
	.I(Ctrl_fsm_data[30]),
	.OEN(IO_sdram_dq_0_6),
	.IO(IO_sdram_dq[30]),
	.O(IO_sdram_dq_in[30])
);
IOBUF IO_sdram_dq_31_iobuf (
	.I(Ctrl_fsm_data[31]),
	.OEN(IO_sdram_dq_0_6),
	.IO(IO_sdram_dq[31]),
	.O(IO_sdram_dq_in[31])
);
LUT3 \u_sdrc_hs_top/O_sdram_ras_n_d_s  (
	.I0(\u_sdrc_hs_top/Sdram_ras_n ),
	.I1(\u_sdrc_hs_top/Sdram_cmd_init [2]),
	.I2(O_sdrc_init_done),
	.F(O_sdram_ras_n)
);
defparam \u_sdrc_hs_top/O_sdram_ras_n_d_s .INIT=8'hAC;
LUT3 \u_sdrc_hs_top/O_sdram_cas_n_d_s  (
	.I0(\u_sdrc_hs_top/Sdram_cmd_init [1]),
	.I1(\u_sdrc_hs_top/Sdram_cas_n ),
	.I2(O_sdrc_init_done),
	.F(O_sdram_cas_n)
);
defparam \u_sdrc_hs_top/O_sdram_cas_n_d_s .INIT=8'hCA;
LUT3 \u_sdrc_hs_top/O_sdram_wen_n_d_s  (
	.I0(\u_sdrc_hs_top/Sdram_cmd_init [0]),
	.I1(\u_sdrc_hs_top/Sdram_wen_n ),
	.I2(O_sdrc_init_done),
	.F(O_sdram_wen_n)
);
defparam \u_sdrc_hs_top/O_sdram_wen_n_d_s .INIT=8'hCA;
LUT3 \u_sdrc_hs_top/O_sdram_addr_d_10_s  (
	.I0(\u_sdrc_hs_top/Sdram_ba_init [1]),
	.I1(\u_sdrc_hs_top/Sdram_addr [10]),
	.I2(O_sdrc_init_done),
	.F(O_sdram_addr[10])
);
defparam \u_sdrc_hs_top/O_sdram_addr_d_10_s .INIT=8'hCA;
LUT3 \u_sdrc_hs_top/O_sdram_addr_d_9_s  (
	.I0(\u_sdrc_hs_top/Sdram_ba_init [1]),
	.I1(\u_sdrc_hs_top/Sdram_addr [9]),
	.I2(O_sdrc_init_done),
	.F(O_sdram_addr[9])
);
defparam \u_sdrc_hs_top/O_sdram_addr_d_9_s .INIT=8'hCA;
LUT3 \u_sdrc_hs_top/O_sdram_addr_d_8_s  (
	.I0(\u_sdrc_hs_top/Sdram_ba_init [1]),
	.I1(\u_sdrc_hs_top/Sdram_addr [8]),
	.I2(O_sdrc_init_done),
	.F(O_sdram_addr[8])
);
defparam \u_sdrc_hs_top/O_sdram_addr_d_8_s .INIT=8'hCA;
LUT3 \u_sdrc_hs_top/O_sdram_addr_d_7_s  (
	.I0(\u_sdrc_hs_top/Sdram_ba_init [1]),
	.I1(\u_sdrc_hs_top/Sdram_addr [7]),
	.I2(O_sdrc_init_done),
	.F(O_sdram_addr[7])
);
defparam \u_sdrc_hs_top/O_sdram_addr_d_7_s .INIT=8'hCA;
LUT3 \u_sdrc_hs_top/O_sdram_addr_d_6_s  (
	.I0(\u_sdrc_hs_top/Sdram_ba_init [1]),
	.I1(\u_sdrc_hs_top/Sdram_addr [6]),
	.I2(O_sdrc_init_done),
	.F(O_sdram_addr[6])
);
defparam \u_sdrc_hs_top/O_sdram_addr_d_6_s .INIT=8'hCA;
LUT3 \u_sdrc_hs_top/O_sdram_addr_d_4_s  (
	.I0(\u_sdrc_hs_top/Sdram_ba_init [1]),
	.I1(\u_sdrc_hs_top/Sdram_addr [4]),
	.I2(O_sdrc_init_done),
	.F(O_sdram_addr[4])
);
defparam \u_sdrc_hs_top/O_sdram_addr_d_4_s .INIT=8'hCA;
LUT3 \u_sdrc_hs_top/O_sdram_addr_d_3_s  (
	.I0(\u_sdrc_hs_top/Sdram_ba_init [1]),
	.I1(\u_sdrc_hs_top/Sdram_addr [3]),
	.I2(O_sdrc_init_done),
	.F(O_sdram_addr[3])
);
defparam \u_sdrc_hs_top/O_sdram_addr_d_3_s .INIT=8'hCA;
LUT3 \u_sdrc_hs_top/O_sdram_addr_d_2_s  (
	.I0(\u_sdrc_hs_top/Sdram_ba_init [1]),
	.I1(\u_sdrc_hs_top/Sdram_addr [2]),
	.I2(O_sdrc_init_done),
	.F(O_sdram_addr[2])
);
defparam \u_sdrc_hs_top/O_sdram_addr_d_2_s .INIT=8'hCA;
LUT3 \u_sdrc_hs_top/O_sdram_addr_d_1_s  (
	.I0(\u_sdrc_hs_top/Sdram_ba_init [1]),
	.I1(\u_sdrc_hs_top/Sdram_addr [1]),
	.I2(O_sdrc_init_done),
	.F(O_sdram_addr[1])
);
defparam \u_sdrc_hs_top/O_sdram_addr_d_1_s .INIT=8'hCA;
LUT3 \u_sdrc_hs_top/O_sdram_addr_d_0_s  (
	.I0(\u_sdrc_hs_top/Sdram_ba_init [1]),
	.I1(\u_sdrc_hs_top/Sdram_addr [0]),
	.I2(O_sdrc_init_done),
	.F(O_sdram_addr[0])
);
defparam \u_sdrc_hs_top/O_sdram_addr_d_0_s .INIT=8'hCA;
LUT3 \u_sdrc_hs_top/O_sdram_ba_d_1_s  (
	.I0(\u_sdrc_hs_top/Sdram_ba_init [1]),
	.I1(\u_sdrc_hs_top/Sdram_ba [1]),
	.I2(O_sdrc_init_done),
	.F(O_sdram_ba[1])
);
defparam \u_sdrc_hs_top/O_sdram_ba_d_1_s .INIT=8'hCA;
LUT3 \u_sdrc_hs_top/O_sdram_ba_d_0_s  (
	.I0(\u_sdrc_hs_top/Sdram_ba_init [1]),
	.I1(\u_sdrc_hs_top/Sdram_ba [0]),
	.I2(O_sdrc_init_done),
	.F(O_sdram_ba[0])
);
defparam \u_sdrc_hs_top/O_sdram_ba_d_0_s .INIT=8'hCA;
LUT3 \u_sdrc_hs_top/n202_s1  (
	.I0(\u_sdrc_hs_top/Cmd_init_state.INIT_STATE_LOAD_MODEREG ),
	.I1(\u_sdrc_hs_top/Cmd_init_state.INIT_STATE_AUTOREFRESH2 ),
	.I2(\u_sdrc_hs_top/Cmd_init_state.INIT_STATE_AUTOREFRESH1 ),
	.F(\u_sdrc_hs_top/n202_5 )
);
defparam \u_sdrc_hs_top/n202_s1 .INIT=8'h01;
LUT2 \u_sdrc_hs_top/n204_s1  (
	.I0(\u_sdrc_hs_top/Cmd_init_state.INIT_STATE_LOAD_MODEREG ),
	.I1(\u_sdrc_hs_top/Cmd_init_state.INIT_STATE_PRECHARGEALL ),
	.F(\u_sdrc_hs_top/n204_5 )
);
defparam \u_sdrc_hs_top/n204_s1 .INIT=4'h1;
LUT4 \u_sdrc_hs_top/n153_s11  (
	.I0(\u_sdrc_hs_top/Cmd_init_state.INIT_STATE_IDLE ),
	.I1(\u_sdrc_hs_top/Init_cnt [15]),
	.I2(\u_sdrc_hs_top/n153_16 ),
	.I3(\u_sdrc_hs_top/Cmd_init_state.INIT_STATE_PRECHARGEALL ),
	.F(\u_sdrc_hs_top/n153_15 )
);
defparam \u_sdrc_hs_top/n153_s11 .INIT=16'h8F88;
LUT4 \u_sdrc_hs_top/n155_s12  (
	.I0(\u_sdrc_hs_top/n155_17 ),
	.I1(\u_sdrc_hs_top/n153_16 ),
	.I2(\u_sdrc_hs_top/Cmd_init_state.INIT_STATE_AUTOREFRESH1 ),
	.I3(\u_sdrc_hs_top/Cmd_init_state.INIT_STATE_PRECHARGE_DELAY ),
	.F(\u_sdrc_hs_top/n155_16 )
);
defparam \u_sdrc_hs_top/n155_s12 .INIT=16'hFA30;
LUT4 \u_sdrc_hs_top/n157_s12  (
	.I0(\u_sdrc_hs_top/n157_17 ),
	.I1(\u_sdrc_hs_top/n153_16 ),
	.I2(\u_sdrc_hs_top/Cmd_init_state.INIT_STATE_AUTOREFRESH2 ),
	.I3(\u_sdrc_hs_top/Cmd_init_state.INIT_STATE_AUTOREFRESH1_DELAY ),
	.F(\u_sdrc_hs_top/n157_16 )
);
defparam \u_sdrc_hs_top/n157_s12 .INIT=16'hFA30;
LUT4 \u_sdrc_hs_top/n159_s12  (
	.I0(\u_sdrc_hs_top/n157_17 ),
	.I1(\u_sdrc_hs_top/n153_16 ),
	.I2(\u_sdrc_hs_top/Cmd_init_state.INIT_STATE_LOAD_MODEREG ),
	.I3(\u_sdrc_hs_top/Cmd_init_state.INIT_STATE_AUTOREFRESH2_DELAY ),
	.F(\u_sdrc_hs_top/n159_16 )
);
defparam \u_sdrc_hs_top/n159_s12 .INIT=16'hFA30;
LUT2 \u_sdrc_hs_top/n161_s11  (
	.I0(\u_sdrc_hs_top/n153_16 ),
	.I1(\u_sdrc_hs_top/Cmd_init_state.INIT_STATE_IDLE ),
	.F(\u_sdrc_hs_top/n161_15 )
);
defparam \u_sdrc_hs_top/n161_s11 .INIT=4'h4;
LUT3 \u_sdrc_hs_top/n163_s12  (
	.I0(\u_sdrc_hs_top/n163_17 ),
	.I1(\u_sdrc_hs_top/Cmd_init_state.INIT_STATE_PRECHARGE_DELAY ),
	.I2(\u_sdrc_hs_top/Cmd_init_state.INIT_STATE_PRECHARGEALL ),
	.F(\u_sdrc_hs_top/n163_16 )
);
defparam \u_sdrc_hs_top/n163_s12 .INIT=8'hF4;
LUT3 \u_sdrc_hs_top/n169_s12  (
	.I0(\u_sdrc_hs_top/n163_17 ),
	.I1(\u_sdrc_hs_top/Cmd_init_state.INIT_STATE_LOAD_MODEREG_DELAY ),
	.I2(\u_sdrc_hs_top/Cmd_init_state.INIT_STATE_LOAD_MODEREG ),
	.F(\u_sdrc_hs_top/n169_16 )
);
defparam \u_sdrc_hs_top/n169_s12 .INIT=8'hF4;
LUT3 \u_sdrc_hs_top/n171_s13  (
	.I0(\u_sdrc_hs_top/Cmd_init_state.INIT_STATE_LOAD_MODEREG_DELAY ),
	.I1(\u_sdrc_hs_top/n155_17 ),
	.I2(\u_sdrc_hs_top/Cmd_init_state.INIT_STATE_INIT_DONE ),
	.F(\u_sdrc_hs_top/n171_17 )
);
defparam \u_sdrc_hs_top/n171_s13 .INIT=8'hF8;
LUT2 \u_sdrc_hs_top/O_sdram_cke_d_s  (
	.I0(\u_sdrc_hs_top/Sdram_cke ),
	.I1(O_sdrc_init_done),
	.F(O_sdram_cke)
);
defparam \u_sdrc_hs_top/O_sdram_cke_d_s .INIT=4'hB;
LUT2 \u_sdrc_hs_top/O_sdram_addr_d_5_s  (
	.I0(\u_sdrc_hs_top/Sdram_addr [5]),
	.I1(O_sdrc_init_done),
	.F(O_sdram_addr[5])
);
defparam \u_sdrc_hs_top/O_sdram_addr_d_5_s .INIT=4'hB;
LUT2 \u_sdrc_hs_top/n65_s0  (
	.I0(\u_sdrc_hs_top/Count_init_delay [0]),
	.I1(\u_sdrc_hs_top/Count_init_delay [1]),
	.F(\u_sdrc_hs_top/n65_4 )
);
defparam \u_sdrc_hs_top/n65_s0 .INIT=4'h6;
LUT3 \u_sdrc_hs_top/n64_s0  (
	.I0(\u_sdrc_hs_top/Count_init_delay [0]),
	.I1(\u_sdrc_hs_top/Count_init_delay [1]),
	.I2(\u_sdrc_hs_top/Count_init_delay [2]),
	.F(\u_sdrc_hs_top/n64_4 )
);
defparam \u_sdrc_hs_top/n64_s0 .INIT=8'h78;
LUT4 \u_sdrc_hs_top/n63_s0  (
	.I0(\u_sdrc_hs_top/Count_init_delay [0]),
	.I1(\u_sdrc_hs_top/Count_init_delay [1]),
	.I2(\u_sdrc_hs_top/Count_init_delay [2]),
	.I3(\u_sdrc_hs_top/Count_init_delay [3]),
	.F(\u_sdrc_hs_top/n63_4 )
);
defparam \u_sdrc_hs_top/n63_s0 .INIT=16'h7F80;
LUT4 \u_sdrc_hs_top/n153_s12  (
	.I0(\u_sdrc_hs_top/Cmd_init_state.INIT_STATE_AUTOREFRESH1_DELAY ),
	.I1(\u_sdrc_hs_top/Cmd_init_state.INIT_STATE_AUTOREFRESH2_DELAY ),
	.I2(\u_sdrc_hs_top/n157_17 ),
	.I3(\u_sdrc_hs_top/n153_17 ),
	.F(\u_sdrc_hs_top/n153_16 )
);
defparam \u_sdrc_hs_top/n153_s12 .INIT=16'hF100;
LUT4 \u_sdrc_hs_top/n155_s13  (
	.I0(\u_sdrc_hs_top/Count_init_delay [0]),
	.I1(\u_sdrc_hs_top/Count_init_delay [2]),
	.I2(\u_sdrc_hs_top/Count_init_delay [3]),
	.I3(\u_sdrc_hs_top/Count_init_delay [1]),
	.F(\u_sdrc_hs_top/n155_17 )
);
defparam \u_sdrc_hs_top/n155_s13 .INIT=16'h0100;
LUT4 \u_sdrc_hs_top/n157_s13  (
	.I0(\u_sdrc_hs_top/Count_init_delay [0]),
	.I1(\u_sdrc_hs_top/Count_init_delay [1]),
	.I2(\u_sdrc_hs_top/Count_init_delay [2]),
	.I3(\u_sdrc_hs_top/Count_init_delay [3]),
	.F(\u_sdrc_hs_top/n157_17 )
);
defparam \u_sdrc_hs_top/n157_s13 .INIT=16'h0100;
LUT4 \u_sdrc_hs_top/n163_s13  (
	.I0(\u_sdrc_hs_top/Cmd_init_state.INIT_STATE_AUTOREFRESH2_DELAY ),
	.I1(\u_sdrc_hs_top/Cmd_init_state.INIT_STATE_AUTOREFRESH1_DELAY ),
	.I2(\u_sdrc_hs_top/n163_18 ),
	.I3(\u_sdrc_hs_top/n155_17 ),
	.F(\u_sdrc_hs_top/n163_17 )
);
defparam \u_sdrc_hs_top/n163_s13 .INIT=16'h0100;
LUT4 \u_sdrc_hs_top/n153_s13  (
	.I0(\u_sdrc_hs_top/Cmd_init_state.INIT_STATE_PRECHARGE_DELAY ),
	.I1(\u_sdrc_hs_top/Cmd_init_state.INIT_STATE_LOAD_MODEREG_DELAY ),
	.I2(\u_sdrc_hs_top/n155_17 ),
	.I3(\u_sdrc_hs_top/n163_18 ),
	.F(\u_sdrc_hs_top/n153_17 )
);
defparam \u_sdrc_hs_top/n153_s13 .INIT=16'h00F1;
LUT2 \u_sdrc_hs_top/n163_s14  (
	.I0(\u_sdrc_hs_top/Init_cnt [15]),
	.I1(\u_sdrc_hs_top/Cmd_init_state.INIT_STATE_IDLE ),
	.F(\u_sdrc_hs_top/n163_18 )
);
defparam \u_sdrc_hs_top/n163_s14 .INIT=4'h4;
LUT4 \u_sdrc_hs_top/n167_s13  (
	.I0(\u_sdrc_hs_top/n153_17 ),
	.I1(\u_sdrc_hs_top/n157_17 ),
	.I2(\u_sdrc_hs_top/Cmd_init_state.INIT_STATE_AUTOREFRESH2_DELAY ),
	.I3(\u_sdrc_hs_top/Cmd_init_state.INIT_STATE_AUTOREFRESH2 ),
	.F(\u_sdrc_hs_top/n167_18 )
);
defparam \u_sdrc_hs_top/n167_s13 .INIT=16'hFF70;
LUT4 \u_sdrc_hs_top/n165_s14  (
	.I0(\u_sdrc_hs_top/n153_17 ),
	.I1(\u_sdrc_hs_top/n157_17 ),
	.I2(\u_sdrc_hs_top/Cmd_init_state.INIT_STATE_AUTOREFRESH1_DELAY ),
	.I3(\u_sdrc_hs_top/Cmd_init_state.INIT_STATE_AUTOREFRESH1 ),
	.F(\u_sdrc_hs_top/n165_19 )
);
defparam \u_sdrc_hs_top/n165_s14 .INIT=16'hFF70;
LUT4 \u_sdrc_hs_top/n200_s2  (
	.I0(\u_sdrc_hs_top/Cmd_init_state.INIT_STATE_PRECHARGEALL ),
	.I1(\u_sdrc_hs_top/Cmd_init_state.INIT_STATE_LOAD_MODEREG ),
	.I2(\u_sdrc_hs_top/Cmd_init_state.INIT_STATE_AUTOREFRESH2 ),
	.I3(\u_sdrc_hs_top/Cmd_init_state.INIT_STATE_AUTOREFRESH1 ),
	.F(\u_sdrc_hs_top/n200_7 )
);
defparam \u_sdrc_hs_top/n200_s2 .INIT=16'h0001;
LUT2 \u_sdrc_hs_top/n27_s3  (
	.I0(\u_sdrc_hs_top/Init_cnt [0]),
	.I1(\u_sdrc_hs_top/Init_cnt [15]),
	.F(\u_sdrc_hs_top/n27_11 )
);
defparam \u_sdrc_hs_top/n27_s3 .INIT=4'h9;
LUT4 \u_sdrc_hs_top/n67_s2  (
	.I0(\u_sdrc_hs_top/Cmd_init_state.INIT_STATE_PRECHARGEALL ),
	.I1(\u_sdrc_hs_top/Cmd_init_state.INIT_STATE_LOAD_MODEREG ),
	.I2(\u_sdrc_hs_top/Cmd_init_state.INIT_STATE_AUTOREFRESH2 ),
	.I3(\u_sdrc_hs_top/Cmd_init_state.INIT_STATE_AUTOREFRESH1 ),
	.F(\u_sdrc_hs_top/n67_6 )
);
defparam \u_sdrc_hs_top/n67_s2 .INIT=16'hFFFE;
DFFCE \u_sdrc_hs_top/Init_cnt_14_s0  (
	.D(\u_sdrc_hs_top/n13_1 ),
	.CLK(I_sdrc_clk),
	.CE(\u_sdrc_hs_top/Init_cnt_14_9 ),
	.CLEAR(\u_sdrc_hs_top/n9_6 ),
	.Q(\u_sdrc_hs_top/Init_cnt [14])
);
defparam \u_sdrc_hs_top/Init_cnt_14_s0 .INIT=1'b0;
DFFCE \u_sdrc_hs_top/Init_cnt_13_s0  (
	.D(\u_sdrc_hs_top/n14_1 ),
	.CLK(I_sdrc_clk),
	.CE(\u_sdrc_hs_top/Init_cnt_14_9 ),
	.CLEAR(\u_sdrc_hs_top/n9_6 ),
	.Q(\u_sdrc_hs_top/Init_cnt [13])
);
defparam \u_sdrc_hs_top/Init_cnt_13_s0 .INIT=1'b0;
DFFCE \u_sdrc_hs_top/Init_cnt_12_s0  (
	.D(\u_sdrc_hs_top/n15_1 ),
	.CLK(I_sdrc_clk),
	.CE(\u_sdrc_hs_top/Init_cnt_14_9 ),
	.CLEAR(\u_sdrc_hs_top/n9_6 ),
	.Q(\u_sdrc_hs_top/Init_cnt [12])
);
defparam \u_sdrc_hs_top/Init_cnt_12_s0 .INIT=1'b0;
DFFCE \u_sdrc_hs_top/Init_cnt_11_s0  (
	.D(\u_sdrc_hs_top/n16_1 ),
	.CLK(I_sdrc_clk),
	.CE(\u_sdrc_hs_top/Init_cnt_14_9 ),
	.CLEAR(\u_sdrc_hs_top/n9_6 ),
	.Q(\u_sdrc_hs_top/Init_cnt [11])
);
defparam \u_sdrc_hs_top/Init_cnt_11_s0 .INIT=1'b0;
DFFCE \u_sdrc_hs_top/Init_cnt_10_s0  (
	.D(\u_sdrc_hs_top/n17_1 ),
	.CLK(I_sdrc_clk),
	.CE(\u_sdrc_hs_top/Init_cnt_14_9 ),
	.CLEAR(\u_sdrc_hs_top/n9_6 ),
	.Q(\u_sdrc_hs_top/Init_cnt [10])
);
defparam \u_sdrc_hs_top/Init_cnt_10_s0 .INIT=1'b0;
DFFCE \u_sdrc_hs_top/Init_cnt_9_s0  (
	.D(\u_sdrc_hs_top/n18_1 ),
	.CLK(I_sdrc_clk),
	.CE(\u_sdrc_hs_top/Init_cnt_14_9 ),
	.CLEAR(\u_sdrc_hs_top/n9_6 ),
	.Q(\u_sdrc_hs_top/Init_cnt [9])
);
defparam \u_sdrc_hs_top/Init_cnt_9_s0 .INIT=1'b0;
DFFCE \u_sdrc_hs_top/Init_cnt_8_s0  (
	.D(\u_sdrc_hs_top/n19_1 ),
	.CLK(I_sdrc_clk),
	.CE(\u_sdrc_hs_top/Init_cnt_14_9 ),
	.CLEAR(\u_sdrc_hs_top/n9_6 ),
	.Q(\u_sdrc_hs_top/Init_cnt [8])
);
defparam \u_sdrc_hs_top/Init_cnt_8_s0 .INIT=1'b0;
DFFCE \u_sdrc_hs_top/Init_cnt_7_s0  (
	.D(\u_sdrc_hs_top/n20_1 ),
	.CLK(I_sdrc_clk),
	.CE(\u_sdrc_hs_top/Init_cnt_14_9 ),
	.CLEAR(\u_sdrc_hs_top/n9_6 ),
	.Q(\u_sdrc_hs_top/Init_cnt [7])
);
defparam \u_sdrc_hs_top/Init_cnt_7_s0 .INIT=1'b0;
DFFCE \u_sdrc_hs_top/Init_cnt_6_s0  (
	.D(\u_sdrc_hs_top/n21_1 ),
	.CLK(I_sdrc_clk),
	.CE(\u_sdrc_hs_top/Init_cnt_14_9 ),
	.CLEAR(\u_sdrc_hs_top/n9_6 ),
	.Q(\u_sdrc_hs_top/Init_cnt [6])
);
defparam \u_sdrc_hs_top/Init_cnt_6_s0 .INIT=1'b0;
DFFCE \u_sdrc_hs_top/Init_cnt_5_s0  (
	.D(\u_sdrc_hs_top/n22_1 ),
	.CLK(I_sdrc_clk),
	.CE(\u_sdrc_hs_top/Init_cnt_14_9 ),
	.CLEAR(\u_sdrc_hs_top/n9_6 ),
	.Q(\u_sdrc_hs_top/Init_cnt [5])
);
defparam \u_sdrc_hs_top/Init_cnt_5_s0 .INIT=1'b0;
DFFCE \u_sdrc_hs_top/Init_cnt_4_s0  (
	.D(\u_sdrc_hs_top/n23_1 ),
	.CLK(I_sdrc_clk),
	.CE(\u_sdrc_hs_top/Init_cnt_14_9 ),
	.CLEAR(\u_sdrc_hs_top/n9_6 ),
	.Q(\u_sdrc_hs_top/Init_cnt [4])
);
defparam \u_sdrc_hs_top/Init_cnt_4_s0 .INIT=1'b0;
DFFCE \u_sdrc_hs_top/Init_cnt_3_s0  (
	.D(\u_sdrc_hs_top/n24_1 ),
	.CLK(I_sdrc_clk),
	.CE(\u_sdrc_hs_top/Init_cnt_14_9 ),
	.CLEAR(\u_sdrc_hs_top/n9_6 ),
	.Q(\u_sdrc_hs_top/Init_cnt [3])
);
defparam \u_sdrc_hs_top/Init_cnt_3_s0 .INIT=1'b0;
DFFCE \u_sdrc_hs_top/Init_cnt_2_s0  (
	.D(\u_sdrc_hs_top/n25_1 ),
	.CLK(I_sdrc_clk),
	.CE(\u_sdrc_hs_top/Init_cnt_14_9 ),
	.CLEAR(\u_sdrc_hs_top/n9_6 ),
	.Q(\u_sdrc_hs_top/Init_cnt [2])
);
defparam \u_sdrc_hs_top/Init_cnt_2_s0 .INIT=1'b0;
DFFCE \u_sdrc_hs_top/Init_cnt_1_s0  (
	.D(\u_sdrc_hs_top/n26_1 ),
	.CLK(I_sdrc_clk),
	.CE(\u_sdrc_hs_top/Init_cnt_14_9 ),
	.CLEAR(\u_sdrc_hs_top/n9_6 ),
	.Q(\u_sdrc_hs_top/Init_cnt [1])
);
defparam \u_sdrc_hs_top/Init_cnt_1_s0 .INIT=1'b0;
DFFR \u_sdrc_hs_top/Count_init_delay_3_s0  (
	.D(\u_sdrc_hs_top/n63_4 ),
	.CLK(I_sdrc_clk),
	.RESET(\u_sdrc_hs_top/n67_6 ),
	.Q(\u_sdrc_hs_top/Count_init_delay [3])
);
defparam \u_sdrc_hs_top/Count_init_delay_3_s0 .INIT=1'b0;
DFFR \u_sdrc_hs_top/Count_init_delay_2_s0  (
	.D(\u_sdrc_hs_top/n64_4 ),
	.CLK(I_sdrc_clk),
	.RESET(\u_sdrc_hs_top/n67_6 ),
	.Q(\u_sdrc_hs_top/Count_init_delay [2])
);
defparam \u_sdrc_hs_top/Count_init_delay_2_s0 .INIT=1'b0;
DFFR \u_sdrc_hs_top/Count_init_delay_1_s0  (
	.D(\u_sdrc_hs_top/n65_4 ),
	.CLK(I_sdrc_clk),
	.RESET(\u_sdrc_hs_top/n67_6 ),
	.Q(\u_sdrc_hs_top/Count_init_delay [1])
);
defparam \u_sdrc_hs_top/Count_init_delay_1_s0 .INIT=1'b0;
DFFR \u_sdrc_hs_top/Count_init_delay_0_s0  (
	.D(\u_sdrc_hs_top/n66_6 ),
	.CLK(I_sdrc_clk),
	.RESET(\u_sdrc_hs_top/n67_6 ),
	.Q(\u_sdrc_hs_top/Count_init_delay [0])
);
defparam \u_sdrc_hs_top/Count_init_delay_0_s0 .INIT=1'b0;
DFFC \u_sdrc_hs_top/Cmd_init_state.INIT_STATE_PRECHARGEALL_s0  (
	.D(\u_sdrc_hs_top/n153_15 ),
	.CLK(I_sdrc_clk),
	.CLEAR(\u_sdrc_hs_top/n9_6 ),
	.Q(\u_sdrc_hs_top/Cmd_init_state.INIT_STATE_PRECHARGEALL )
);
defparam \u_sdrc_hs_top/Cmd_init_state.INIT_STATE_PRECHARGEALL_s0 .INIT=1'b0;
DFFC \u_sdrc_hs_top/Cmd_init_state.INIT_STATE_AUTOREFRESH1_s0  (
	.D(\u_sdrc_hs_top/n155_16 ),
	.CLK(I_sdrc_clk),
	.CLEAR(\u_sdrc_hs_top/n9_6 ),
	.Q(\u_sdrc_hs_top/Cmd_init_state.INIT_STATE_AUTOREFRESH1 )
);
defparam \u_sdrc_hs_top/Cmd_init_state.INIT_STATE_AUTOREFRESH1_s0 .INIT=1'b0;
DFFC \u_sdrc_hs_top/Cmd_init_state.INIT_STATE_AUTOREFRESH2_s0  (
	.D(\u_sdrc_hs_top/n157_16 ),
	.CLK(I_sdrc_clk),
	.CLEAR(\u_sdrc_hs_top/n9_6 ),
	.Q(\u_sdrc_hs_top/Cmd_init_state.INIT_STATE_AUTOREFRESH2 )
);
defparam \u_sdrc_hs_top/Cmd_init_state.INIT_STATE_AUTOREFRESH2_s0 .INIT=1'b0;
DFFC \u_sdrc_hs_top/Cmd_init_state.INIT_STATE_LOAD_MODEREG_s0  (
	.D(\u_sdrc_hs_top/n159_16 ),
	.CLK(I_sdrc_clk),
	.CLEAR(\u_sdrc_hs_top/n9_6 ),
	.Q(\u_sdrc_hs_top/Cmd_init_state.INIT_STATE_LOAD_MODEREG )
);
defparam \u_sdrc_hs_top/Cmd_init_state.INIT_STATE_LOAD_MODEREG_s0 .INIT=1'b0;
DFFC \u_sdrc_hs_top/Cmd_init_state.INIT_STATE_PRECHARGE_DELAY_s0  (
	.D(\u_sdrc_hs_top/n163_16 ),
	.CLK(I_sdrc_clk),
	.CLEAR(\u_sdrc_hs_top/n9_6 ),
	.Q(\u_sdrc_hs_top/Cmd_init_state.INIT_STATE_PRECHARGE_DELAY )
);
defparam \u_sdrc_hs_top/Cmd_init_state.INIT_STATE_PRECHARGE_DELAY_s0 .INIT=1'b0;
DFFC \u_sdrc_hs_top/Cmd_init_state.INIT_STATE_AUTOREFRESH1_DELAY_s0  (
	.D(\u_sdrc_hs_top/n165_19 ),
	.CLK(I_sdrc_clk),
	.CLEAR(\u_sdrc_hs_top/n9_6 ),
	.Q(\u_sdrc_hs_top/Cmd_init_state.INIT_STATE_AUTOREFRESH1_DELAY )
);
defparam \u_sdrc_hs_top/Cmd_init_state.INIT_STATE_AUTOREFRESH1_DELAY_s0 .INIT=1'b0;
DFFC \u_sdrc_hs_top/Cmd_init_state.INIT_STATE_AUTOREFRESH2_DELAY_s0  (
	.D(\u_sdrc_hs_top/n167_18 ),
	.CLK(I_sdrc_clk),
	.CLEAR(\u_sdrc_hs_top/n9_6 ),
	.Q(\u_sdrc_hs_top/Cmd_init_state.INIT_STATE_AUTOREFRESH2_DELAY )
);
defparam \u_sdrc_hs_top/Cmd_init_state.INIT_STATE_AUTOREFRESH2_DELAY_s0 .INIT=1'b0;
DFFC \u_sdrc_hs_top/Cmd_init_state.INIT_STATE_LOAD_MODEREG_DELAY_s0  (
	.D(\u_sdrc_hs_top/n169_16 ),
	.CLK(I_sdrc_clk),
	.CLEAR(\u_sdrc_hs_top/n9_6 ),
	.Q(\u_sdrc_hs_top/Cmd_init_state.INIT_STATE_LOAD_MODEREG_DELAY )
);
defparam \u_sdrc_hs_top/Cmd_init_state.INIT_STATE_LOAD_MODEREG_DELAY_s0 .INIT=1'b0;
DFFC \u_sdrc_hs_top/Cmd_init_state.INIT_STATE_INIT_DONE_s0  (
	.D(\u_sdrc_hs_top/n171_17 ),
	.CLK(I_sdrc_clk),
	.CLEAR(\u_sdrc_hs_top/n9_6 ),
	.Q(\u_sdrc_hs_top/Cmd_init_state.INIT_STATE_INIT_DONE )
);
defparam \u_sdrc_hs_top/Cmd_init_state.INIT_STATE_INIT_DONE_s0 .INIT=1'b0;
DFFC \u_sdrc_hs_top/Init_finish_s0  (
	.D(\u_sdrc_hs_top/Cmd_init_state.INIT_STATE_INIT_DONE ),
	.CLK(I_sdrc_clk),
	.CLEAR(\u_sdrc_hs_top/n9_6 ),
	.Q(O_sdrc_init_done)
);
defparam \u_sdrc_hs_top/Init_finish_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/Sdram_cmd_init_2_s0  (
	.D(\u_sdrc_hs_top/n200_7 ),
	.CLK(I_sdrc_clk),
	.Q(\u_sdrc_hs_top/Sdram_cmd_init [2])
);
defparam \u_sdrc_hs_top/Sdram_cmd_init_2_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/Sdram_cmd_init_1_s0  (
	.D(\u_sdrc_hs_top/n202_5 ),
	.CLK(I_sdrc_clk),
	.Q(\u_sdrc_hs_top/Sdram_cmd_init [1])
);
defparam \u_sdrc_hs_top/Sdram_cmd_init_1_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/Sdram_cmd_init_0_s0  (
	.D(\u_sdrc_hs_top/n204_5 ),
	.CLK(I_sdrc_clk),
	.Q(\u_sdrc_hs_top/Sdram_cmd_init [0])
);
defparam \u_sdrc_hs_top/Sdram_cmd_init_0_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/Sdram_ba_init_1_s0  (
	.D(\u_sdrc_hs_top/n205_6 ),
	.CLK(I_sdrc_clk),
	.Q(\u_sdrc_hs_top/Sdram_ba_init [1])
);
defparam \u_sdrc_hs_top/Sdram_ba_init_1_s0 .INIT=1'b0;
DFFP \u_sdrc_hs_top/Cmd_init_state.INIT_STATE_IDLE_s0  (
	.D(\u_sdrc_hs_top/n161_15 ),
	.CLK(I_sdrc_clk),
	.PRESET(\u_sdrc_hs_top/n9_6 ),
	.Q(\u_sdrc_hs_top/Cmd_init_state.INIT_STATE_IDLE )
);
defparam \u_sdrc_hs_top/Cmd_init_state.INIT_STATE_IDLE_s0 .INIT=1'b1;
DFFCE \u_sdrc_hs_top/Init_cnt_15_s1  (
	.D(VCC),
	.CLK(I_sdrc_clk),
	.CE(\u_sdrc_hs_top/n12_1 ),
	.CLEAR(\u_sdrc_hs_top/n9_6 ),
	.Q(\u_sdrc_hs_top/Init_cnt [15])
);
defparam \u_sdrc_hs_top/Init_cnt_15_s1 .INIT=1'b0;
DFFC \u_sdrc_hs_top/Init_cnt_0_s2  (
	.D(\u_sdrc_hs_top/n27_11 ),
	.CLK(I_sdrc_clk),
	.CLEAR(\u_sdrc_hs_top/n9_6 ),
	.Q(\u_sdrc_hs_top/Init_cnt [0])
);
defparam \u_sdrc_hs_top/Init_cnt_0_s2 .INIT=1'b0;
ODDR \u_sdrc_hs_top/U_ODDR_clk  (
	.D0(VCC),
	.D1(GND),
	.CLK(I_sdram_clk),
	.TX(VCC),
	.Q0(O_sdram_clk),
	.Q1(\u_sdrc_hs_top/U_ODDR_clk_1_Q1 )
);
defparam \u_sdrc_hs_top/U_ODDR_clk .INIT=1'b0;
defparam \u_sdrc_hs_top/U_ODDR_clk .TXCLK_POL=1'b0;
ALU \u_sdrc_hs_top/n26_s  (
	.I0(\u_sdrc_hs_top/Init_cnt [1]),
	.I1(\u_sdrc_hs_top/Init_cnt [0]),
	.I3(GND),
	.CIN(GND),
	.COUT(\u_sdrc_hs_top/n26_2 ),
	.SUM(\u_sdrc_hs_top/n26_1 )
);
defparam \u_sdrc_hs_top/n26_s .ALU_MODE=0;
ALU \u_sdrc_hs_top/n25_s  (
	.I0(GND),
	.I1(\u_sdrc_hs_top/Init_cnt [2]),
	.I3(GND),
	.CIN(\u_sdrc_hs_top/n26_2 ),
	.COUT(\u_sdrc_hs_top/n25_2 ),
	.SUM(\u_sdrc_hs_top/n25_1 )
);
defparam \u_sdrc_hs_top/n25_s .ALU_MODE=0;
ALU \u_sdrc_hs_top/n24_s  (
	.I0(GND),
	.I1(\u_sdrc_hs_top/Init_cnt [3]),
	.I3(GND),
	.CIN(\u_sdrc_hs_top/n25_2 ),
	.COUT(\u_sdrc_hs_top/n24_2 ),
	.SUM(\u_sdrc_hs_top/n24_1 )
);
defparam \u_sdrc_hs_top/n24_s .ALU_MODE=0;
ALU \u_sdrc_hs_top/n23_s  (
	.I0(GND),
	.I1(\u_sdrc_hs_top/Init_cnt [4]),
	.I3(GND),
	.CIN(\u_sdrc_hs_top/n24_2 ),
	.COUT(\u_sdrc_hs_top/n23_2 ),
	.SUM(\u_sdrc_hs_top/n23_1 )
);
defparam \u_sdrc_hs_top/n23_s .ALU_MODE=0;
ALU \u_sdrc_hs_top/n22_s  (
	.I0(GND),
	.I1(\u_sdrc_hs_top/Init_cnt [5]),
	.I3(GND),
	.CIN(\u_sdrc_hs_top/n23_2 ),
	.COUT(\u_sdrc_hs_top/n22_2 ),
	.SUM(\u_sdrc_hs_top/n22_1 )
);
defparam \u_sdrc_hs_top/n22_s .ALU_MODE=0;
ALU \u_sdrc_hs_top/n21_s  (
	.I0(GND),
	.I1(\u_sdrc_hs_top/Init_cnt [6]),
	.I3(GND),
	.CIN(\u_sdrc_hs_top/n22_2 ),
	.COUT(\u_sdrc_hs_top/n21_2 ),
	.SUM(\u_sdrc_hs_top/n21_1 )
);
defparam \u_sdrc_hs_top/n21_s .ALU_MODE=0;
ALU \u_sdrc_hs_top/n20_s  (
	.I0(GND),
	.I1(\u_sdrc_hs_top/Init_cnt [7]),
	.I3(GND),
	.CIN(\u_sdrc_hs_top/n21_2 ),
	.COUT(\u_sdrc_hs_top/n20_2 ),
	.SUM(\u_sdrc_hs_top/n20_1 )
);
defparam \u_sdrc_hs_top/n20_s .ALU_MODE=0;
ALU \u_sdrc_hs_top/n19_s  (
	.I0(GND),
	.I1(\u_sdrc_hs_top/Init_cnt [8]),
	.I3(GND),
	.CIN(\u_sdrc_hs_top/n20_2 ),
	.COUT(\u_sdrc_hs_top/n19_2 ),
	.SUM(\u_sdrc_hs_top/n19_1 )
);
defparam \u_sdrc_hs_top/n19_s .ALU_MODE=0;
ALU \u_sdrc_hs_top/n18_s  (
	.I0(GND),
	.I1(\u_sdrc_hs_top/Init_cnt [9]),
	.I3(GND),
	.CIN(\u_sdrc_hs_top/n19_2 ),
	.COUT(\u_sdrc_hs_top/n18_2 ),
	.SUM(\u_sdrc_hs_top/n18_1 )
);
defparam \u_sdrc_hs_top/n18_s .ALU_MODE=0;
ALU \u_sdrc_hs_top/n17_s  (
	.I0(GND),
	.I1(\u_sdrc_hs_top/Init_cnt [10]),
	.I3(GND),
	.CIN(\u_sdrc_hs_top/n18_2 ),
	.COUT(\u_sdrc_hs_top/n17_2 ),
	.SUM(\u_sdrc_hs_top/n17_1 )
);
defparam \u_sdrc_hs_top/n17_s .ALU_MODE=0;
ALU \u_sdrc_hs_top/n16_s  (
	.I0(GND),
	.I1(\u_sdrc_hs_top/Init_cnt [11]),
	.I3(GND),
	.CIN(\u_sdrc_hs_top/n17_2 ),
	.COUT(\u_sdrc_hs_top/n16_2 ),
	.SUM(\u_sdrc_hs_top/n16_1 )
);
defparam \u_sdrc_hs_top/n16_s .ALU_MODE=0;
ALU \u_sdrc_hs_top/n15_s  (
	.I0(GND),
	.I1(\u_sdrc_hs_top/Init_cnt [12]),
	.I3(GND),
	.CIN(\u_sdrc_hs_top/n16_2 ),
	.COUT(\u_sdrc_hs_top/n15_2 ),
	.SUM(\u_sdrc_hs_top/n15_1 )
);
defparam \u_sdrc_hs_top/n15_s .ALU_MODE=0;
ALU \u_sdrc_hs_top/n14_s  (
	.I0(GND),
	.I1(\u_sdrc_hs_top/Init_cnt [13]),
	.I3(GND),
	.CIN(\u_sdrc_hs_top/n15_2 ),
	.COUT(\u_sdrc_hs_top/n14_2 ),
	.SUM(\u_sdrc_hs_top/n14_1 )
);
defparam \u_sdrc_hs_top/n14_s .ALU_MODE=0;
ALU \u_sdrc_hs_top/n13_s  (
	.I0(GND),
	.I1(\u_sdrc_hs_top/Init_cnt [14]),
	.I3(GND),
	.CIN(\u_sdrc_hs_top/n14_2 ),
	.COUT(\u_sdrc_hs_top/n13_2 ),
	.SUM(\u_sdrc_hs_top/n13_1 )
);
defparam \u_sdrc_hs_top/n13_s .ALU_MODE=0;
ALU \u_sdrc_hs_top/n12_s  (
	.I0(GND),
	.I1(\u_sdrc_hs_top/Init_cnt [15]),
	.I3(GND),
	.CIN(\u_sdrc_hs_top/n13_2 ),
	.COUT(\u_sdrc_hs_top/n12_0_COUT ),
	.SUM(\u_sdrc_hs_top/n12_1 )
);
defparam \u_sdrc_hs_top/n12_s .ALU_MODE=0;
INV \u_sdrc_hs_top/n9_s2  (
	.I(I_sdrc_rst_n),
	.O(\u_sdrc_hs_top/n9_6 )
);
LUT1 \u_sdrc_hs_top/n205_s2  (
	.I0(\u_sdrc_hs_top/Cmd_init_state.INIT_STATE_LOAD_MODEREG ),
	.F(\u_sdrc_hs_top/n205_6 )
);
defparam \u_sdrc_hs_top/n205_s2 .INIT=2'h1;
LUT1 \u_sdrc_hs_top/n66_s2  (
	.I0(\u_sdrc_hs_top/Count_init_delay [0]),
	.F(\u_sdrc_hs_top/n66_6 )
);
defparam \u_sdrc_hs_top/n66_s2 .INIT=2'h1;
INV \u_sdrc_hs_top/Init_cnt_14_s4  (
	.I(\u_sdrc_hs_top/Init_cnt [15]),
	.O(\u_sdrc_hs_top/Init_cnt_14_9 )
);
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/n179_s0  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n179_4 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n179_5 ),
	.I2(I_sdrc_cmd_en),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n179_3 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n179_s0 .INIT=8'hCA;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n180_s0  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n180_10 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd [6]),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n180_8 ),
	.I3(I_sdrc_cmd_en),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n180_3 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n180_s0 .INIT=16'hAA3C;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n181_s0  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n181_8 ),
	.I1(I_sdrc_addr[5]),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n181_5 ),
	.I3(I_sdrc_cmd_en),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n181_3 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n181_s0 .INIT=16'h3CAA;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n182_s0  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n182_4 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd [4]),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n182_5 ),
	.I3(I_sdrc_cmd_en),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n182_3 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n182_s0 .INIT=16'hAA3C;
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/n183_s0  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n183_7 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n183_5 ),
	.I2(I_sdrc_cmd_en),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n183_3 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n183_s0 .INIT=8'hCA;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n184_s0  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n184_4 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd [2]),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n184_5 ),
	.I3(I_sdrc_cmd_en),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n184_3 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n184_s0 .INIT=16'hAA3C;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n185_s0  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n185_4 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd [0]),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd [1]),
	.I3(I_sdrc_cmd_en),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n185_3 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n185_s0 .INIT=16'hAA3C;
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/n186_s0  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd [0]),
	.I1(I_sdrc_addr[0]),
	.I2(I_sdrc_cmd_en),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n186_3 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n186_s0 .INIT=8'h35;
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_wr_data_valid_s3  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_WRITE_WITHOUT_AUTOPRE ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_wr_data_valid_9 ),
	.I2(I_sdrc_cmd_en),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_wr_data_valid_8 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_wr_data_valid_s3 .INIT=8'hF8;
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/n80_s25  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n606_17 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_DATAIN2ACTIVE ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n80_32 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n80_29 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n80_s25 .INIT=8'hBF;
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/n590_s27  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n590_32 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_DATAIN2ACTIVE ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n590_33 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n590_31 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n590_s27 .INIT=8'hF4;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n592_s27  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n592_40 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n592_33 ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n592_38 ),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/n592_35 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n592_31 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n592_s27 .INIT=16'hFF07;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n997_s12  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_wr_data_valid_9 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_WRITE_WITHOUT_AUTOPRE ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n997_17 ),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/n997_18 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n997_16 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n997_s12 .INIT=16'hF8FF;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1003_s12  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n1003_17 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_IDLE ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n997_17 ),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/n1003_18 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1003_16 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1003_s12 .INIT=16'hF4FF;
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/n580_s28  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n590_32 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_AUTOREFRESH_DELAY ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n580_36 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n580_32 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n580_s28 .INIT=8'hF4;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n582_s27  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_32 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_33 ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_34 ),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_35 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_31 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n582_s27 .INIT=16'hEFFF;
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/n584_s28  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n590_32 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_ACTIVE2RW_DELAY ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n584_33 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n584_32 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n584_s28 .INIT=8'hF4;
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/n586_s27  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n586_32 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_READ_WITHOUT_AUTOPRE ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n586_33 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n586_31 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n586_s27 .INIT=8'hF4;
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/n588_s27  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n586_32 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_WRITE_WITHOUT_AUTOPRE ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n588_32 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n588_31 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n588_s27 .INIT=8'hF4;
LUT2 \u_sdrc_hs_top/u_sdrc_control_fsm/n594_s27  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n590_32 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_INIT ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n594_31 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n594_s27 .INIT=4'h4;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n596_s29  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n590_32 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_POWER_DOWN ),
	.I2(I_sdram_power_down),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_IDLE ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n596_33 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n596_s29 .INIT=16'hF444;
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/n598_s29  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n592_40 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_SELFREFRESH ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n598_34 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n598_33 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n598_s29 .INIT=8'hF4;
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/n602_s28  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n590_32 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_SELFREFRESH_WAIT ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_SELFREFRESH ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n602_32 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n602_s28 .INIT=8'hF4;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n604_s27  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n590_32 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_SELFREFRESH_EXIT ),
	.I2(I_sdram_selfrefresh),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_SELFREFRESH_WAIT ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n604_31 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n604_s27 .INIT=16'h4F44;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1000_s13  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_wr_data_valid_9 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd_7_9 ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n1000_18 ),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/n1000_19 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1000_17 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1000_s13 .INIT=16'hF2FF;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1005_s14  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n1005_19 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_IDLE ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n1005_20 ),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/n1005_21 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1005_18 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1005_s14 .INIT=16'h8FFF;
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/n1007_s14  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n1007_19 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n1005_20 ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n1007_20 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1007_18 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1007_s14 .INIT=8'hBF;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1009_s14  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n1009_24 ),
	.I1(\u_sdrc_hs_top/Sdram_addr [10]),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n1009_20 ),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/n1005_20 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1009_18 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1009_s14 .INIT=16'hF4FF;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1011_s14  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n1009_24 ),
	.I1(\u_sdrc_hs_top/Sdram_addr [9]),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n1011_19 ),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/n1005_20 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1011_18 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1011_s14 .INIT=16'hF4FF;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1013_s14  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n1009_24 ),
	.I1(\u_sdrc_hs_top/Sdram_addr [8]),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n1013_19 ),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/n1005_20 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1013_18 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1013_s14 .INIT=16'hF4FF;
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/n1015_s14  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n1015_19 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n1005_20 ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n1015_20 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1015_18 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1015_s14 .INIT=8'hBF;
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/n1017_s14  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n1017_19 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n1005_20 ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n1017_20 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1017_18 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1017_s14 .INIT=8'hBF;
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/n1019_s14  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n1019_19 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n1005_20 ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n1019_20 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1019_18 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1019_s14 .INIT=8'hBF;
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/n1021_s14  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n1021_19 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n1005_20 ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n1021_20 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1021_18 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1021_s14 .INIT=8'hBF;
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/n1023_s14  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n1023_19 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n1005_20 ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n1023_20 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1023_18 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1023_s14 .INIT=8'hBF;
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/n1025_s14  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n1025_19 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n1005_20 ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n1025_20 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1025_18 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1025_s14 .INIT=8'hBF;
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/n1027_s14  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n1027_19 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n1005_20 ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n1027_20 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1027_18 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1027_s14 .INIT=8'hBF;
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/n1029_s14  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n1029_19 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n1005_20 ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n1029_20 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1029_18 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1029_s14 .INIT=8'hBF;
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/n80_s26  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n80_33 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_34 ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n80_34 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n80_31 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n80_s26 .INIT=8'hBF;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n606_s9  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num [7]),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n606_19 ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd_7_9 ),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num [8]),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n606_14 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n606_s9 .INIT=16'h0708;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n618_s8  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num [0]),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num [1]),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd_7_9 ),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num [2]),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n618_12 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n618_s8 .INIT=16'h0708;
LUT2 \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_cke_s5  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_cke_8 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_DATAIN2ACTIVE ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_cke_7 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_cke_s5 .INIT=4'hB;
LUT2 \u_sdrc_hs_top/u_sdrc_control_fsm/n86_s0  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay [0]),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay [1]),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n86_4 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n86_s0 .INIT=4'h6;
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/n85_s0  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay [0]),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay [1]),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay [2]),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n85_4 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n85_s0 .INIT=8'h78;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n84_s0  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay [0]),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay [1]),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay [2]),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay [3]),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n84_4 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n84_s0 .INIT=16'h7F80;
LUT2 \u_sdrc_hs_top/u_sdrc_control_fsm/n100_s0  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay2 [0]),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay2 [1]),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n100_4 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n100_s0 .INIT=4'h6;
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/n99_s0  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay2 [0]),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay2 [1]),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay2 [2]),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n99_4 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n99_s0 .INIT=8'h78;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n98_s0  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay2 [0]),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay2 [1]),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay2 [2]),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay2 [3]),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n98_4 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n98_s0 .INIT=16'h7F80;
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/n179_s1  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd [6]),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n180_8 ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd [7]),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n179_4 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n179_s1 .INIT=8'h78;
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/n179_s2  (
	.I0(I_sdrc_addr[6]),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n179_8 ),
	.I2(I_sdrc_addr[7]),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n179_5 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n179_s2 .INIT=8'h78;
LUT2 \u_sdrc_hs_top/u_sdrc_control_fsm/n181_s2  (
	.I0(I_sdrc_addr[4]),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n181_6 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n181_5 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n181_s2 .INIT=4'h8;
LUT2 \u_sdrc_hs_top/u_sdrc_control_fsm/n182_s1  (
	.I0(I_sdrc_addr[4]),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n181_6 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n182_4 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n182_s1 .INIT=4'h6;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n182_s2  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd [0]),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd [1]),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd [2]),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd [3]),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n182_5 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n182_s2 .INIT=16'h8000;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n183_s2  (
	.I0(I_sdrc_addr[0]),
	.I1(I_sdrc_addr[2]),
	.I2(I_sdrc_addr[1]),
	.I3(I_sdrc_addr[3]),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n183_5 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n183_s2 .INIT=16'h7F80;
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/n184_s1  (
	.I0(I_sdrc_addr[0]),
	.I1(I_sdrc_addr[1]),
	.I2(I_sdrc_addr[2]),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n184_4 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n184_s1 .INIT=8'h78;
LUT2 \u_sdrc_hs_top/u_sdrc_control_fsm/n184_s2  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd [0]),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd [1]),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n184_5 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n184_s2 .INIT=4'h8;
LUT2 \u_sdrc_hs_top/u_sdrc_control_fsm/n185_s1  (
	.I0(I_sdrc_addr[0]),
	.I1(I_sdrc_addr[1]),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n185_4 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n185_s1 .INIT=4'h6;
LUT2 \u_sdrc_hs_top/u_sdrc_control_fsm/n993_s1  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_DATAIN2ACTIVE ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n993_5 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n993_4 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n993_s1 .INIT=4'h4;
LUT2 \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd_7_s4  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_WRITE_WITHOUT_AUTOPRE ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_READ_WITHOUT_AUTOPRE ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd_7_9 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd_7_s4 .INIT=4'h1;
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_wr_data_valid_s4  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_wr_data_valid_10 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_wr_data_valid_11 ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_wr_data_valid_12 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_wr_data_valid_9 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_wr_data_valid_s4 .INIT=8'h80;
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/n80_s27  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_PRECHARGE_DELAY ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_ACTIVE2RW_DELAY ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_AUTOREFRESH_DELAY ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n80_32 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n80_s27 .INIT=8'h01;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n590_s28  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_wr_data_valid_9 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd_7_9 ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_32 ),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/n590_34 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n590_32 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n590_s28 .INIT=16'h0E00;
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/n590_s29  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Precharge_flag ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_wr_data_valid_9 ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_WRITE_WITHOUT_AUTOPRE ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n590_33 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n590_s29 .INIT=8'h80;
LUT2 \u_sdrc_hs_top/u_sdrc_control_fsm/n592_s29  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_DATAIN2ACTIVE ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_32 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n592_33 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n592_s29 .INIT=4'h1;
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/n592_s31  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_READ_WITHOUT_AUTOPRE ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Precharge_flag ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_wr_data_valid_9 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n592_35 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n592_s31 .INIT=8'h80;
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/n997_s13  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_wr_data_valid_9 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Precharge_flag ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_READ_WITHOUT_AUTOPRE ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n997_17 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n997_s13 .INIT=8'h70;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n997_s14  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_cke_7 ),
	.I1(\u_sdrc_hs_top/Sdram_wen_n ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n997_19 ),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/n997_20 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n997_18 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n997_s14 .INIT=16'h0B00;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1003_s13  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n1003_19 ),
	.I1(\u_sdrc_hs_top/Sdram_ras_n ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n1003_20 ),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/n1003_25 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1003_17 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1003_s13 .INIT=16'hB303;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1003_s14  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_cke_7 ),
	.I1(\u_sdrc_hs_top/Sdram_ras_n ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_WRITE_WITHOUT_AUTOPRE ),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/n1003_22 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1003_18 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1003_s14 .INIT=16'h0B00;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n582_s28  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n1003_19 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_36 ),
	.I2(I_sdrc_cmd_en),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_54 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_32 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n582_s28 .INIT=16'h1F00;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n582_s29  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd_7_9 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_wr_data_valid_9 ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_38 ),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_IDLE ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_33 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n582_s29 .INIT=16'h1F00;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n582_s30  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd_7_9 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Precharge_flag ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_wr_data_valid_9 ),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_39 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_34 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n582_s30 .INIT=16'h00EF;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n582_s31  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_40 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_AUTOREFRESH_DELAY ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_41 ),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_42 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_35 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n582_s31 .INIT=16'h7000;
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/n584_s29  (
	.I0(I_sdrc_cmd[1]),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_54 ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n584_36 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n584_33 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n584_s29 .INIT=8'h80;
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/n586_s28  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_32 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_wr_data_valid_9 ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n590_34 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n586_32 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n586_s28 .INIT=8'h40;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n586_s29  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n586_34 ),
	.I1(I_sdrc_cmd[0]),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n759_6 ),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/n580_38 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n586_33 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n586_s29 .INIT=16'h4000;
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/n588_s28  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n586_34 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_54 ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n759_8 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n588_32 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n588_s28 .INIT=8'h40;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n598_s30  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n584_36 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_SELFREFRESH ),
	.I2(I_sdram_selfrefresh),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/n598_35 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n598_34 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n598_s30 .INIT=16'hF400;
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/n1000_s14  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n1000_20 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n1000_21 ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_IDLE ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1000_18 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1000_s14 .INIT=8'hD0;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1000_s15  (
	.I0(\u_sdrc_hs_top/Sdram_cas_n ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_cke_8 ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_DATAIN2ACTIVE ),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/n1003_22 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1000_19 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1000_s15 .INIT=16'h1F00;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1005_s15  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n1005_22 ),
	.I1(I_sdrc_cmd_en),
	.I2(\u_sdrc_hs_top/Sdram_ba [1]),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/n1003_20 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1005_19 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1005_s15 .INIT=16'hBBF0;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1005_s16  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_wr_data_valid_9 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd_7_9 ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n592_36 ),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/n997_20 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1005_20 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1005_s16 .INIT=16'h0D00;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1005_s17  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd_7_9 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_bk_wrd [1]),
	.I2(\u_sdrc_hs_top/Sdram_ba [1]),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_DATAIN2ACTIVE ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1005_21 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1005_s17 .INIT=16'h0BBB;
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/n1007_s15  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n1007_21 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n1007_22 ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_IDLE ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1007_19 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1007_s15 .INIT=8'h10;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1007_s16  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd_7_9 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_bk_wrd [0]),
	.I2(\u_sdrc_hs_top/Sdram_ba [0]),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_DATAIN2ACTIVE ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1007_20 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1007_s16 .INIT=16'h0BBB;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1009_s16  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n759_6 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n1009_21 ),
	.I2(I_sdrc_cmd_en),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_54 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1009_20 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1009_s16 .INIT=16'h4F00;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1011_s15  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n759_6 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n1011_20 ),
	.I2(I_sdrc_cmd_en),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_54 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1011_19 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1011_s15 .INIT=16'h4F00;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1013_s15  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n759_6 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n1013_20 ),
	.I2(I_sdrc_cmd_en),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_54 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1013_19 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1013_s15 .INIT=16'h4F00;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1015_s15  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n1015_21 ),
	.I1(\u_sdrc_hs_top/Sdram_addr [7]),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n1003_20 ),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_IDLE ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1015_19 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1015_s15 .INIT=16'h5C00;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1015_s16  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd_7_9 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd [7]),
	.I2(\u_sdrc_hs_top/Sdram_addr [7]),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_DATAIN2ACTIVE ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1015_20 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1015_s16 .INIT=16'h0BBB;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1017_s15  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n1017_21 ),
	.I1(\u_sdrc_hs_top/Sdram_addr [6]),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n1003_20 ),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_IDLE ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1017_19 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1017_s15 .INIT=16'h5C00;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1017_s16  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd_7_9 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd [6]),
	.I2(\u_sdrc_hs_top/Sdram_addr [6]),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_DATAIN2ACTIVE ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1017_20 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1017_s16 .INIT=16'h0BBB;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1019_s15  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n1019_21 ),
	.I1(\u_sdrc_hs_top/Sdram_addr [5]),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n1003_20 ),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_IDLE ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1019_19 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1019_s15 .INIT=16'h5C00;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1019_s16  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd_7_9 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd [5]),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_DATAIN2ACTIVE ),
	.I3(\u_sdrc_hs_top/Sdram_addr [5]),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1019_20 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1019_s16 .INIT=16'h0BBB;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1021_s15  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n1021_21 ),
	.I1(\u_sdrc_hs_top/Sdram_addr [4]),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n1003_20 ),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_IDLE ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1021_19 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1021_s15 .INIT=16'h5C00;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1021_s16  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd_7_9 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd [4]),
	.I2(\u_sdrc_hs_top/Sdram_addr [4]),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_DATAIN2ACTIVE ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1021_20 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1021_s16 .INIT=16'h0BBB;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1023_s15  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n1023_21 ),
	.I1(\u_sdrc_hs_top/Sdram_addr [3]),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n1003_20 ),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_IDLE ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1023_19 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1023_s15 .INIT=16'h5C00;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1023_s16  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd_7_9 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd [3]),
	.I2(\u_sdrc_hs_top/Sdram_addr [3]),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_DATAIN2ACTIVE ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1023_20 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1023_s16 .INIT=16'h0BBB;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1025_s15  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n1025_21 ),
	.I1(\u_sdrc_hs_top/Sdram_addr [2]),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n1003_20 ),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_IDLE ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1025_19 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1025_s15 .INIT=16'h5C00;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1025_s16  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd_7_9 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd [2]),
	.I2(\u_sdrc_hs_top/Sdram_addr [2]),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_DATAIN2ACTIVE ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1025_20 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1025_s16 .INIT=16'h0BBB;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1027_s15  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n1027_21 ),
	.I1(\u_sdrc_hs_top/Sdram_addr [1]),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n1003_20 ),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_IDLE ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1027_19 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1027_s15 .INIT=16'h5C00;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1027_s16  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd_7_9 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd [1]),
	.I2(\u_sdrc_hs_top/Sdram_addr [1]),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_DATAIN2ACTIVE ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1027_20 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1027_s16 .INIT=16'h0BBB;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1029_s15  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n1029_21 ),
	.I1(\u_sdrc_hs_top/Sdram_addr [0]),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n1003_20 ),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_IDLE ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1029_19 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1029_s15 .INIT=16'h5C00;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1029_s16  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd_7_9 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd [0]),
	.I2(\u_sdrc_hs_top/Sdram_addr [0]),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_DATAIN2ACTIVE ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1029_20 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1029_s16 .INIT=16'h0BBB;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n80_s28  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n586_34 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n759_6 ),
	.I2(O_sdrc_cmd_ack),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/n580_38 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n80_33 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n80_s28 .INIT=16'hF800;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n80_s29  (
	.I0(O_sdrc_cmd_ack),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_40 ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_AUTOREFRESH_DELAY ),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/n80_35 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n80_34 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n80_s29 .INIT=16'h001F;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n614_s9  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num [0]),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num [1]),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num [2]),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num [3]),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n614_13 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n614_s9 .INIT=16'h8000;
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/n616_s9  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num [0]),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num [1]),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num [2]),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n616_13 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n616_s9 .INIT=8'h80;
LUT2 \u_sdrc_hs_top/u_sdrc_control_fsm/n759_s2  (
	.I0(I_sdrc_cmd[1]),
	.I1(I_sdrc_cmd[2]),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n759_6 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n759_s2 .INIT=4'h4;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_cke_s6  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay2 [1]),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay2 [2]),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay2 [3]),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay2 [0]),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_cke_8 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_cke_s6 .INIT=16'h0100;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n181_s3  (
	.I0(I_sdrc_addr[0]),
	.I1(I_sdrc_addr[3]),
	.I2(I_sdrc_addr[2]),
	.I3(I_sdrc_addr[1]),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n181_6 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n181_s3 .INIT=16'h8000;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n993_s2  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_POWER_DOWN ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_SELFREFRESH ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_SELFREFRESH_WAIT ),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_SELFREFRESH_EXIT ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n993_5 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n993_s2 .INIT=16'h0001;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_wr_data_valid_s5  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num [3]),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Sdrc_wrd_len [3]),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num [4]),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/Sdrc_wrd_len [4]),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_wr_data_valid_10 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_wr_data_valid_s5 .INIT=16'h9009;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_wr_data_valid_s6  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num [0]),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Sdrc_wrd_len [0]),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num [2]),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/Sdrc_wrd_len [2]),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_wr_data_valid_11 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_wr_data_valid_s6 .INIT=16'h9009;
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_wr_data_valid_s7  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num [8]),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_wr_data_valid_13 ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_wr_data_valid_14 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_wr_data_valid_12 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_wr_data_valid_s7 .INIT=8'h40;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n590_s30  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_40 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_AUTOREFRESH_DELAY ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_38 ),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/n590_35 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n590_34 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n590_s30 .INIT=16'hB000;
LUT2 \u_sdrc_hs_top/u_sdrc_control_fsm/n592_s32  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_DATAIN2ACTIVE ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_cke_8 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n592_36 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n592_s32 .INIT=4'h8;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n997_s15  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n759_8 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n1003_20 ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n997_24 ),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_IDLE ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n997_19 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n997_s15 .INIT=16'h0700;
LUT2 \u_sdrc_hs_top/u_sdrc_control_fsm/n997_s16  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Reset_cmd_count ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n993_5 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n997_20 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n997_s16 .INIT=4'h8;
LUT2 \u_sdrc_hs_top/u_sdrc_control_fsm/n1003_s15  (
	.I0(I_sdrc_cmd[2]),
	.I1(I_sdrc_cmd[0]),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1003_19 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1003_s15 .INIT=4'h4;
LUT2 \u_sdrc_hs_top/u_sdrc_control_fsm/n1003_s16  (
	.I0(I_sdram_power_down),
	.I1(I_sdram_selfrefresh),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1003_20 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1003_s16 .INIT=4'h1;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1003_s18  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_SELFREFRESH_EXIT ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Reset_cmd_count ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_SELFREFRESH ),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/n1003_23 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1003_22 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1003_s18 .INIT=16'hFE00;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n582_s32  (
	.I0(I_sdrc_precharge_ctrl),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_43 ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_44 ),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/n759_6 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_36 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n582_s32 .INIT=16'hBF00;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n582_s34  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_cke_8 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_DATAIN2ACTIVE ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_45 ),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_46 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_38 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n582_s34 .INIT=16'h0B00;
LUT2 \u_sdrc_hs_top/u_sdrc_control_fsm/n582_s35  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_ACTIVE2RW_DELAY ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_47 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_39 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n582_s35 .INIT=4'h8;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n582_s36  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay [3]),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay [1]),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay [2]),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay [0]),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_40 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n582_s36 .INIT=16'h4000;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n582_s37  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd_7_9 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n993_4 ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_IDLE ),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_52 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_41 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n582_s37 .INIT=16'hF70F;
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/n582_s38  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_49 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_PRECHARGE_DELAY ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_50 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_42 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n582_s38 .INIT=8'h70;
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/n586_s30  (
	.I0(I_sdrc_precharge_ctrl),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_44 ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_43 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n586_34 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n586_s30 .INIT=8'h40;
LUT2 \u_sdrc_hs_top/u_sdrc_control_fsm/n598_s31  (
	.I0(I_sdram_power_down),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_IDLE ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n598_35 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n598_s31 .INIT=4'h4;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1000_s16  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n1000_22 ),
	.I1(\u_sdrc_hs_top/Sdram_cas_n ),
	.I2(I_sdrc_cmd_en),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/n1003_20 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1000_20 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1000_s16 .INIT=16'h7033;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1000_s17  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n1003_20 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n1003_19 ),
	.I2(\u_sdrc_hs_top/Sdram_cas_n ),
	.I3(I_sdrc_cmd[1]),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1000_21 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1000_s17 .INIT=16'hF800;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1005_s18  (
	.I0(I_sdrc_addr[20]),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n1005_23 ),
	.I2(\u_sdrc_hs_top/Sdram_ba [1]),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/n1005_24 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1005_22 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1005_s18 .INIT=16'hE0EE;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1007_s17  (
	.I0(I_sdrc_addr[19]),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n1005_23 ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n1003_20 ),
	.I3(I_sdrc_cmd_en),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1007_21 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1007_s17 .INIT=16'h1000;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1007_s18  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n1005_24 ),
	.I1(I_sdrc_cmd_en),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n1003_20 ),
	.I3(\u_sdrc_hs_top/Sdram_ba [0]),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1007_22 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1007_s18 .INIT=16'h008F;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1009_s17  (
	.I0(I_sdrc_addr[18]),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n1009_22 ),
	.I2(\u_sdrc_hs_top/Sdram_addr [10]),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/n1003_19 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1009_21 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1009_s17 .INIT=16'hBBB0;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1011_s16  (
	.I0(I_sdrc_addr[17]),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n1009_22 ),
	.I2(\u_sdrc_hs_top/Sdram_addr [9]),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/n1003_19 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1011_20 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1011_s16 .INIT=16'hBBB0;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1013_s16  (
	.I0(I_sdrc_addr[16]),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n1009_22 ),
	.I2(\u_sdrc_hs_top/Sdram_addr [8]),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/n1003_19 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1013_20 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1013_s16 .INIT=16'hBBB0;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1015_s17  (
	.I0(I_sdrc_addr[7]),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n759_6 ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n1015_22 ),
	.I3(I_sdrc_cmd_en),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1015_21 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1015_s17 .INIT=16'h4F00;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1017_s17  (
	.I0(I_sdrc_addr[6]),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n759_6 ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n1017_22 ),
	.I3(I_sdrc_cmd_en),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1017_21 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1017_s17 .INIT=16'h4F00;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1019_s17  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n1019_22 ),
	.I1(I_sdrc_cmd[1]),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n1019_23 ),
	.I3(I_sdrc_cmd_en),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1019_21 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1019_s17 .INIT=16'h4F00;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1021_s17  (
	.I0(I_sdrc_addr[4]),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n759_6 ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n1021_22 ),
	.I3(I_sdrc_cmd_en),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1021_21 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1021_s17 .INIT=16'h4F00;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1023_s17  (
	.I0(I_sdrc_addr[3]),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n759_6 ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n1023_22 ),
	.I3(I_sdrc_cmd_en),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1023_21 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1023_s17 .INIT=16'h4F00;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1025_s17  (
	.I0(I_sdrc_addr[2]),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n759_6 ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n1025_22 ),
	.I3(I_sdrc_cmd_en),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1025_21 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1025_s17 .INIT=16'h4F00;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1027_s17  (
	.I0(I_sdrc_addr[1]),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n759_6 ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n1027_22 ),
	.I3(I_sdrc_cmd_en),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1027_21 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1027_s17 .INIT=16'h4F00;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1029_s17  (
	.I0(I_sdrc_addr[0]),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n759_6 ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n1029_22 ),
	.I3(I_sdrc_cmd_en),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1029_21 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1029_s17 .INIT=16'h4F00;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n80_s30  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_49 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n80_38 ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_PRECHARGE_DELAY ),
	.I3(O_sdrc_cmd_ack),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n80_35 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n80_s30 .INIT=16'hF3A0;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_wr_data_valid_s8  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num [1]),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Sdrc_wrd_len [1]),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num [5]),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/Sdrc_wrd_len [5]),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_wr_data_valid_13 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_wr_data_valid_s8 .INIT=16'h9009;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_wr_data_valid_s9  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num [6]),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Sdrc_wrd_len [6]),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num [7]),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/Sdrc_wrd_len [7]),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_wr_data_valid_14 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_wr_data_valid_s9 .INIT=16'h9009;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n590_s31  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_47 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_ACTIVE2RW_DELAY ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_49 ),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_PRECHARGE_DELAY ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n590_35 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n590_s31 .INIT=16'hB0BB;
LUT2 \u_sdrc_hs_top/u_sdrc_control_fsm/n1003_s19  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_POWER_DOWN ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_SELFREFRESH_WAIT ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1003_23 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1003_s19 .INIT=4'h1;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n582_s39  (
	.I0(I_sdrc_data_len[0]),
	.I1(I_sdrc_data_len[1]),
	.I2(I_sdrc_data_len[2]),
	.I3(I_sdrc_data_len[3]),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_43 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n582_s39 .INIT=16'h0001;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n582_s40  (
	.I0(I_sdrc_data_len[4]),
	.I1(I_sdrc_data_len[5]),
	.I2(I_sdrc_data_len[6]),
	.I3(I_sdrc_data_len[7]),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_44 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n582_s40 .INIT=16'h0001;
LUT2 \u_sdrc_hs_top/u_sdrc_control_fsm/n582_s41  (
	.I0(I_sdram_power_down),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_POWER_DOWN ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_45 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n582_s41 .INIT=4'h8;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n582_s42  (
	.I0(I_sdram_selfrefresh),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_SELFREFRESH_WAIT ),
	.I2(O_sdrc_init_done),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_INIT ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_46 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n582_s42 .INIT=16'h7077;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n582_s43  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay [0]),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay [2]),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay [3]),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay [1]),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_47 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n582_s43 .INIT=16'h0100;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n582_s45  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay [1]),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay [2]),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay [3]),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay [0]),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_49 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n582_s45 .INIT=16'h0100;
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/n582_s46  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_INIT ),
	.I1(O_sdrc_init_done),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_SELFREFRESH_EXIT ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_50 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n582_s46 .INIT=8'h07;
LUT2 \u_sdrc_hs_top/u_sdrc_control_fsm/n1000_s18  (
	.I0(I_sdrc_cmd[0]),
	.I1(I_sdrc_cmd[2]),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1000_22 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1000_s18 .INIT=4'h1;
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/n1005_s19  (
	.I0(I_sdrc_cmd[0]),
	.I1(I_sdrc_cmd[2]),
	.I2(I_sdrc_cmd[1]),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1005_23 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1005_s19 .INIT=8'hD3;
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/n1005_s20  (
	.I0(I_sdrc_cmd[1]),
	.I1(I_sdrc_cmd[0]),
	.I2(I_sdrc_cmd[2]),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1005_24 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1005_s20 .INIT=8'hA3;
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/n1009_s18  (
	.I0(I_sdrc_cmd[2]),
	.I1(I_sdrc_cmd[1]),
	.I2(I_sdrc_cmd[0]),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1009_22 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1009_s18 .INIT=8'h40;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1015_s18  (
	.I0(I_sdrc_addr[15]),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n1009_22 ),
	.I2(\u_sdrc_hs_top/Sdram_addr [7]),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/n1005_24 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1015_22 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1015_s18 .INIT=16'hB0BB;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1017_s18  (
	.I0(I_sdrc_addr[14]),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n1009_22 ),
	.I2(\u_sdrc_hs_top/Sdram_addr [6]),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/n1005_24 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1017_22 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1017_s18 .INIT=16'hB0BB;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1019_s18  (
	.I0(I_sdrc_addr[13]),
	.I1(I_sdrc_cmd[0]),
	.I2(\u_sdrc_hs_top/Sdram_addr [5]),
	.I3(I_sdrc_cmd[2]),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1019_22 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1019_s18 .INIT=16'hF0BB;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1019_s19  (
	.I0(I_sdrc_addr[5]),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n759_6 ),
	.I2(\u_sdrc_hs_top/Sdram_addr [5]),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/n1000_22 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1019_23 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1019_s19 .INIT=16'hB0BB;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1021_s18  (
	.I0(I_sdrc_addr[12]),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n1009_22 ),
	.I2(\u_sdrc_hs_top/Sdram_addr [4]),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/n1005_24 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1021_22 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1021_s18 .INIT=16'hB0BB;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1023_s18  (
	.I0(I_sdrc_addr[11]),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n1009_22 ),
	.I2(\u_sdrc_hs_top/Sdram_addr [3]),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/n1005_24 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1023_22 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1023_s18 .INIT=16'hB0BB;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1025_s18  (
	.I0(I_sdrc_addr[10]),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n1009_22 ),
	.I2(\u_sdrc_hs_top/Sdram_addr [2]),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/n1005_24 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1025_22 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1025_s18 .INIT=16'hB0BB;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1027_s18  (
	.I0(I_sdrc_addr[9]),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n1009_22 ),
	.I2(\u_sdrc_hs_top/Sdram_addr [1]),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/n1005_24 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1027_22 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1027_s18 .INIT=16'hB0BB;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1029_s18  (
	.I0(I_sdrc_addr[8]),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n1009_22 ),
	.I2(\u_sdrc_hs_top/Sdram_addr [0]),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/n1005_24 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1029_22 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1029_s18 .INIT=16'hB0BB;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n997_s18  (
	.I0(I_sdrc_cmd[1]),
	.I1(I_sdrc_cmd[2]),
	.I2(I_sdrc_cmd[0]),
	.I3(I_sdrc_cmd_en),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n997_22 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n997_s18 .INIT=16'h8F00;
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/n181_s4  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd [5]),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd [4]),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n182_5 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n181_8 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n181_s4 .INIT=8'h6A;
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/n180_s4  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd [5]),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd [4]),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n182_5 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n180_8 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n180_s4 .INIT=8'h80;
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/n179_s4  (
	.I0(I_sdrc_addr[5]),
	.I1(I_sdrc_addr[4]),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n181_6 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n179_8 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n179_s4 .INIT=8'h80;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n183_s3  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd [2]),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd [0]),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd [1]),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd [3]),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n183_7 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n183_s3 .INIT=16'h7F80;
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/n592_s33  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_PRECHARGE_DELAY ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_DATAIN2ACTIVE ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_cke_8 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n592_38 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n592_s33 .INIT=8'h15;
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/n610_s10  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num [5]),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num [4]),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/n614_13 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n610_15 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n610_s10 .INIT=8'h80;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n612_s10  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd_7_9 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num [5]),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num [4]),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/n614_13 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n612_15 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n612_s10 .INIT=16'h1444;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n582_s47  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_INIT ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_PRECHARGE_DELAY ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_ACTIVE2RW_DELAY ),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_AUTOREFRESH_DELAY ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_52 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n582_s47 .INIT=16'h0001;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n993_s3  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_SELFREFRESH_EXIT ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/n606_17 ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_DATAIN2ACTIVE ),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/n993_5 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n993_7 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n993_s3 .INIT=16'hEFEE;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n584_s31  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_36 ),
	.I1(I_sdrc_cmd[2]),
	.I2(I_sdrc_cmd[0]),
	.I3(I_sdrc_cmd_en),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n584_36 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n584_s31 .INIT=16'hBA00;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n580_s31  (
	.I0(I_sdrc_cmd[1]),
	.I1(I_sdrc_cmd[2]),
	.I2(I_sdrc_cmd[0]),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/n580_38 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n580_36 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n580_s31 .INIT=16'h1000;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/Reset_cmd_count_s1  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_DATAIN2ACTIVE ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_WRITE_WITHOUT_AUTOPRE ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_READ_WITHOUT_AUTOPRE ),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_IDLE ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/Reset_cmd_count )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Reset_cmd_count_s1 .INIT=16'hFFFE;
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/n1003_s20  (
	.I0(I_sdrc_cmd[1]),
	.I1(I_sdrc_cmd[2]),
	.I2(I_sdrc_cmd_en),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1003_25 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1003_s20 .INIT=8'hB0;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n759_s3  (
	.I0(I_sdrc_cmd[0]),
	.I1(I_sdrc_cmd_en),
	.I2(I_sdrc_cmd[1]),
	.I3(I_sdrc_cmd[2]),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n759_8 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n759_s3 .INIT=16'h0400;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n997_s19  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/n997_22 ),
	.I1(I_sdram_power_down),
	.I2(I_sdram_selfrefresh),
	.I3(\u_sdrc_hs_top/Sdram_wen_n ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n997_24 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n997_s19 .INIT=16'h00FE;
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/n582_s48  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_IDLE ),
	.I1(I_sdram_power_down),
	.I2(I_sdram_selfrefresh),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_54 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n582_s48 .INIT=8'h02;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n1009_s19  (
	.I0(I_sdram_power_down),
	.I1(I_sdram_selfrefresh),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_IDLE ),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_DATAIN2ACTIVE ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n1009_24 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n1009_s19 .INIT=16'h001F;
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/n80_s32  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_ACTIVE2RW_DELAY ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_WRITE_WITHOUT_AUTOPRE ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_READ_WITHOUT_AUTOPRE ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n80_38 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n80_s32 .INIT=8'h01;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n592_s34  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_wr_data_valid_9 ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_WRITE_WITHOUT_AUTOPRE ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_READ_WITHOUT_AUTOPRE ),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/n590_34 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n592_40 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n592_s34 .INIT=16'hAB00;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n620_s9  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_WRITE_WITHOUT_AUTOPRE ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_READ_WITHOUT_AUTOPRE ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num [0]),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num [1]),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n620_14 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n620_s9 .INIT=16'h0EE0;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n616_s10  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_WRITE_WITHOUT_AUTOPRE ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_READ_WITHOUT_AUTOPRE ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num [3]),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/n616_13 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n616_15 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n616_s10 .INIT=16'h0EE0;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n614_s10  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_WRITE_WITHOUT_AUTOPRE ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_READ_WITHOUT_AUTOPRE ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num [4]),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/n614_13 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n614_15 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n614_s10 .INIT=16'h0EE0;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n610_s11  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_WRITE_WITHOUT_AUTOPRE ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_READ_WITHOUT_AUTOPRE ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num [6]),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/n610_15 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n610_17 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n610_s11 .INIT=16'h0EE0;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n608_s9  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_WRITE_WITHOUT_AUTOPRE ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_READ_WITHOUT_AUTOPRE ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num [7]),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/n606_19 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n608_14 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n608_s9 .INIT=16'h0EE0;
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd_7_s5  (
	.I0(I_sdrc_cmd_en),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_WRITE_WITHOUT_AUTOPRE ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_READ_WITHOUT_AUTOPRE ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd_7_11 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd_7_s5 .INIT=8'hFE;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n622_s11  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num [0]),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_WRITE_WITHOUT_AUTOPRE ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_READ_WITHOUT_AUTOPRE ),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_IDLE ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n622_17 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n622_s11 .INIT=16'h5456;
LUT3 \u_sdrc_hs_top/u_sdrc_control_fsm/n606_s11  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_WRITE_WITHOUT_AUTOPRE ),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_READ_WITHOUT_AUTOPRE ),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_IDLE ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n606_17 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n606_s11 .INIT=8'hFE;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n180_s5  (
	.I0(I_sdrc_addr[6]),
	.I1(I_sdrc_addr[5]),
	.I2(I_sdrc_addr[4]),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/n181_6 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n180_10 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n180_s5 .INIT=16'h6AAA;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n606_s12  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num [6]),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num [5]),
	.I2(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num [4]),
	.I3(\u_sdrc_hs_top/u_sdrc_control_fsm/n614_13 ),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n606_19 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n606_s12 .INIT=16'h8000;
LUT4 \u_sdrc_hs_top/u_sdrc_control_fsm/n580_s32  (
	.I0(I_sdrc_cmd_en),
	.I1(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_IDLE ),
	.I2(I_sdram_power_down),
	.I3(I_sdram_selfrefresh),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n580_38 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n580_s32 .INIT=16'h0008;
DFFR \u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay_3_s0  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n84_4 ),
	.CLK(I_sdrc_clk),
	.RESET(\u_sdrc_hs_top/u_sdrc_control_fsm/Reset_cmd_count ),
	.Q(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay [3])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay_3_s0 .INIT=1'b0;
DFFR \u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay_2_s0  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n85_4 ),
	.CLK(I_sdrc_clk),
	.RESET(\u_sdrc_hs_top/u_sdrc_control_fsm/Reset_cmd_count ),
	.Q(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay [2])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay_2_s0 .INIT=1'b0;
DFFR \u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay_1_s0  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n86_4 ),
	.CLK(I_sdrc_clk),
	.RESET(\u_sdrc_hs_top/u_sdrc_control_fsm/Reset_cmd_count ),
	.Q(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay [1])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay_1_s0 .INIT=1'b0;
DFFS \u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay_0_s0  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n87_6 ),
	.CLK(I_sdrc_clk),
	.SET(\u_sdrc_hs_top/u_sdrc_control_fsm/Reset_cmd_count ),
	.Q(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay [0])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay_0_s0 .INIT=1'b1;
DFFR \u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay2_3_s0  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n98_4 ),
	.CLK(I_sdrc_clk),
	.RESET(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_WRITE_WITHOUT_AUTOPRE ),
	.Q(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay2 [3])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay2_3_s0 .INIT=1'b0;
DFFR \u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay2_2_s0  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n99_4 ),
	.CLK(I_sdrc_clk),
	.RESET(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_WRITE_WITHOUT_AUTOPRE ),
	.Q(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay2 [2])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay2_2_s0 .INIT=1'b0;
DFFR \u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay2_1_s0  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n100_4 ),
	.CLK(I_sdrc_clk),
	.RESET(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_WRITE_WITHOUT_AUTOPRE ),
	.Q(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay2 [1])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay2_1_s0 .INIT=1'b0;
DFFS \u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay2_0_s0  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n101_6 ),
	.CLK(I_sdrc_clk),
	.SET(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_WRITE_WITHOUT_AUTOPRE ),
	.Q(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay2 [0])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay2_0_s0 .INIT=1'b1;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_31_s0  (
	.D(I_sdrc_data[31]),
	.CLK(I_sdrc_clk),
	.Q(Ctrl_fsm_data[31])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_31_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_30_s0  (
	.D(I_sdrc_data[30]),
	.CLK(I_sdrc_clk),
	.Q(Ctrl_fsm_data[30])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_30_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_29_s0  (
	.D(I_sdrc_data[29]),
	.CLK(I_sdrc_clk),
	.Q(Ctrl_fsm_data[29])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_29_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_28_s0  (
	.D(I_sdrc_data[28]),
	.CLK(I_sdrc_clk),
	.Q(Ctrl_fsm_data[28])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_28_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_27_s0  (
	.D(I_sdrc_data[27]),
	.CLK(I_sdrc_clk),
	.Q(Ctrl_fsm_data[27])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_27_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_26_s0  (
	.D(I_sdrc_data[26]),
	.CLK(I_sdrc_clk),
	.Q(Ctrl_fsm_data[26])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_26_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_25_s0  (
	.D(I_sdrc_data[25]),
	.CLK(I_sdrc_clk),
	.Q(Ctrl_fsm_data[25])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_25_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_24_s0  (
	.D(I_sdrc_data[24]),
	.CLK(I_sdrc_clk),
	.Q(Ctrl_fsm_data[24])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_24_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_23_s0  (
	.D(I_sdrc_data[23]),
	.CLK(I_sdrc_clk),
	.Q(Ctrl_fsm_data[23])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_23_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_22_s0  (
	.D(I_sdrc_data[22]),
	.CLK(I_sdrc_clk),
	.Q(Ctrl_fsm_data[22])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_22_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_21_s0  (
	.D(I_sdrc_data[21]),
	.CLK(I_sdrc_clk),
	.Q(Ctrl_fsm_data[21])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_21_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_20_s0  (
	.D(I_sdrc_data[20]),
	.CLK(I_sdrc_clk),
	.Q(Ctrl_fsm_data[20])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_20_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_19_s0  (
	.D(I_sdrc_data[19]),
	.CLK(I_sdrc_clk),
	.Q(Ctrl_fsm_data[19])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_19_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_18_s0  (
	.D(I_sdrc_data[18]),
	.CLK(I_sdrc_clk),
	.Q(Ctrl_fsm_data[18])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_18_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_17_s0  (
	.D(I_sdrc_data[17]),
	.CLK(I_sdrc_clk),
	.Q(Ctrl_fsm_data[17])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_17_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_16_s0  (
	.D(I_sdrc_data[16]),
	.CLK(I_sdrc_clk),
	.Q(Ctrl_fsm_data[16])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_16_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_15_s0  (
	.D(I_sdrc_data[15]),
	.CLK(I_sdrc_clk),
	.Q(Ctrl_fsm_data[15])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_15_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_14_s0  (
	.D(I_sdrc_data[14]),
	.CLK(I_sdrc_clk),
	.Q(Ctrl_fsm_data[14])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_14_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_13_s0  (
	.D(I_sdrc_data[13]),
	.CLK(I_sdrc_clk),
	.Q(Ctrl_fsm_data[13])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_13_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_12_s0  (
	.D(I_sdrc_data[12]),
	.CLK(I_sdrc_clk),
	.Q(Ctrl_fsm_data[12])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_12_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_11_s0  (
	.D(I_sdrc_data[11]),
	.CLK(I_sdrc_clk),
	.Q(Ctrl_fsm_data[11])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_11_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_10_s0  (
	.D(I_sdrc_data[10]),
	.CLK(I_sdrc_clk),
	.Q(Ctrl_fsm_data[10])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_10_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_9_s0  (
	.D(I_sdrc_data[9]),
	.CLK(I_sdrc_clk),
	.Q(Ctrl_fsm_data[9])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_9_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_8_s0  (
	.D(I_sdrc_data[8]),
	.CLK(I_sdrc_clk),
	.Q(Ctrl_fsm_data[8])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_8_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_7_s0  (
	.D(I_sdrc_data[7]),
	.CLK(I_sdrc_clk),
	.Q(Ctrl_fsm_data[7])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_7_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_6_s0  (
	.D(I_sdrc_data[6]),
	.CLK(I_sdrc_clk),
	.Q(Ctrl_fsm_data[6])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_6_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_5_s0  (
	.D(I_sdrc_data[5]),
	.CLK(I_sdrc_clk),
	.Q(Ctrl_fsm_data[5])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_5_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_4_s0  (
	.D(I_sdrc_data[4]),
	.CLK(I_sdrc_clk),
	.Q(Ctrl_fsm_data[4])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_4_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_3_s0  (
	.D(I_sdrc_data[3]),
	.CLK(I_sdrc_clk),
	.Q(Ctrl_fsm_data[3])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_3_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_2_s0  (
	.D(I_sdrc_data[2]),
	.CLK(I_sdrc_clk),
	.Q(Ctrl_fsm_data[2])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_2_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_1_s0  (
	.D(I_sdrc_data[1]),
	.CLK(I_sdrc_clk),
	.Q(Ctrl_fsm_data[1])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_1_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_0_s0  (
	.D(I_sdrc_data[0]),
	.CLK(I_sdrc_clk),
	.Q(Ctrl_fsm_data[0])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_data_0_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_dqm_3_s0  (
	.D(I_sdrc_dqm[3]),
	.CLK(I_sdrc_clk),
	.Q(O_sdram_dqm[3])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_dqm_3_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_dqm_2_s0  (
	.D(I_sdrc_dqm[2]),
	.CLK(I_sdrc_clk),
	.Q(O_sdram_dqm[2])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_dqm_2_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_dqm_1_s0  (
	.D(I_sdrc_dqm[1]),
	.CLK(I_sdrc_clk),
	.Q(O_sdram_dqm[1])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_dqm_1_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_dqm_0_s0  (
	.D(I_sdrc_dqm[0]),
	.CLK(I_sdrc_clk),
	.Q(O_sdram_dqm[0])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_dqm_0_s0 .INIT=1'b0;
DFFE \u_sdrc_hs_top/u_sdrc_control_fsm/Precharge_flag_s0  (
	.D(I_sdrc_precharge_ctrl),
	.CLK(I_sdrc_clk),
	.CE(I_sdrc_cmd_en),
	.Q(\u_sdrc_hs_top/u_sdrc_control_fsm/Precharge_flag )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Precharge_flag_s0 .INIT=1'b0;
DFFE \u_sdrc_hs_top/u_sdrc_control_fsm/Sdrc_wrd_len_7_s0  (
	.D(I_sdrc_data_len[7]),
	.CLK(I_sdrc_clk),
	.CE(I_sdrc_cmd_en),
	.Q(\u_sdrc_hs_top/u_sdrc_control_fsm/Sdrc_wrd_len [7])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Sdrc_wrd_len_7_s0 .INIT=1'b0;
DFFE \u_sdrc_hs_top/u_sdrc_control_fsm/Sdrc_wrd_len_6_s0  (
	.D(I_sdrc_data_len[6]),
	.CLK(I_sdrc_clk),
	.CE(I_sdrc_cmd_en),
	.Q(\u_sdrc_hs_top/u_sdrc_control_fsm/Sdrc_wrd_len [6])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Sdrc_wrd_len_6_s0 .INIT=1'b0;
DFFE \u_sdrc_hs_top/u_sdrc_control_fsm/Sdrc_wrd_len_5_s0  (
	.D(I_sdrc_data_len[5]),
	.CLK(I_sdrc_clk),
	.CE(I_sdrc_cmd_en),
	.Q(\u_sdrc_hs_top/u_sdrc_control_fsm/Sdrc_wrd_len [5])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Sdrc_wrd_len_5_s0 .INIT=1'b0;
DFFE \u_sdrc_hs_top/u_sdrc_control_fsm/Sdrc_wrd_len_4_s0  (
	.D(I_sdrc_data_len[4]),
	.CLK(I_sdrc_clk),
	.CE(I_sdrc_cmd_en),
	.Q(\u_sdrc_hs_top/u_sdrc_control_fsm/Sdrc_wrd_len [4])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Sdrc_wrd_len_4_s0 .INIT=1'b0;
DFFE \u_sdrc_hs_top/u_sdrc_control_fsm/Sdrc_wrd_len_3_s0  (
	.D(I_sdrc_data_len[3]),
	.CLK(I_sdrc_clk),
	.CE(I_sdrc_cmd_en),
	.Q(\u_sdrc_hs_top/u_sdrc_control_fsm/Sdrc_wrd_len [3])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Sdrc_wrd_len_3_s0 .INIT=1'b0;
DFFE \u_sdrc_hs_top/u_sdrc_control_fsm/Sdrc_wrd_len_2_s0  (
	.D(I_sdrc_data_len[2]),
	.CLK(I_sdrc_clk),
	.CE(I_sdrc_cmd_en),
	.Q(\u_sdrc_hs_top/u_sdrc_control_fsm/Sdrc_wrd_len [2])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Sdrc_wrd_len_2_s0 .INIT=1'b0;
DFFE \u_sdrc_hs_top/u_sdrc_control_fsm/Sdrc_wrd_len_1_s0  (
	.D(I_sdrc_data_len[1]),
	.CLK(I_sdrc_clk),
	.CE(I_sdrc_cmd_en),
	.Q(\u_sdrc_hs_top/u_sdrc_control_fsm/Sdrc_wrd_len [1])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Sdrc_wrd_len_1_s0 .INIT=1'b0;
DFFE \u_sdrc_hs_top/u_sdrc_control_fsm/Sdrc_wrd_len_0_s0  (
	.D(I_sdrc_data_len[0]),
	.CLK(I_sdrc_clk),
	.CE(I_sdrc_cmd_en),
	.Q(\u_sdrc_hs_top/u_sdrc_control_fsm/Sdrc_wrd_len [0])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Sdrc_wrd_len_0_s0 .INIT=1'b0;
DFFE \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_bk_wrd_1_s0  (
	.D(I_sdrc_addr[20]),
	.CLK(I_sdrc_clk),
	.CE(I_sdrc_cmd_en),
	.Q(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_bk_wrd [1])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_bk_wrd_1_s0 .INIT=1'b0;
DFFE \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_bk_wrd_0_s0  (
	.D(I_sdrc_addr[19]),
	.CLK(I_sdrc_clk),
	.CE(I_sdrc_cmd_en),
	.Q(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_bk_wrd [0])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_bk_wrd_0_s0 .INIT=1'b0;
DFFC \u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_AUTOREFRESH_DELAY_s0  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n580_32 ),
	.CLK(I_sdrc_clk),
	.CLEAR(\u_sdrc_hs_top/n9_6 ),
	.Q(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_AUTOREFRESH_DELAY )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_AUTOREFRESH_DELAY_s0 .INIT=1'b0;
DFFC \u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_IDLE_s0  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n582_31 ),
	.CLK(I_sdrc_clk),
	.CLEAR(\u_sdrc_hs_top/n9_6 ),
	.Q(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_IDLE )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_IDLE_s0 .INIT=1'b0;
DFFC \u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_ACTIVE2RW_DELAY_s0  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n584_32 ),
	.CLK(I_sdrc_clk),
	.CLEAR(\u_sdrc_hs_top/n9_6 ),
	.Q(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_ACTIVE2RW_DELAY )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_ACTIVE2RW_DELAY_s0 .INIT=1'b0;
DFFC \u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_READ_WITHOUT_AUTOPRE_s0  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n586_31 ),
	.CLK(I_sdrc_clk),
	.CLEAR(\u_sdrc_hs_top/n9_6 ),
	.Q(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_READ_WITHOUT_AUTOPRE )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_READ_WITHOUT_AUTOPRE_s0 .INIT=1'b0;
DFFC \u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_WRITE_WITHOUT_AUTOPRE_s0  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n588_31 ),
	.CLK(I_sdrc_clk),
	.CLEAR(\u_sdrc_hs_top/n9_6 ),
	.Q(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_WRITE_WITHOUT_AUTOPRE )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_WRITE_WITHOUT_AUTOPRE_s0 .INIT=1'b0;
DFFC \u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_DATAIN2ACTIVE_s0  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n590_31 ),
	.CLK(I_sdrc_clk),
	.CLEAR(\u_sdrc_hs_top/n9_6 ),
	.Q(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_DATAIN2ACTIVE )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_DATAIN2ACTIVE_s0 .INIT=1'b0;
DFFC \u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_PRECHARGE_DELAY_s0  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n592_31 ),
	.CLK(I_sdrc_clk),
	.CLEAR(\u_sdrc_hs_top/n9_6 ),
	.Q(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_PRECHARGE_DELAY )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_PRECHARGE_DELAY_s0 .INIT=1'b0;
DFFP \u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_INIT_s0  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n594_31 ),
	.CLK(I_sdrc_clk),
	.PRESET(\u_sdrc_hs_top/n9_6 ),
	.Q(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_INIT )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_INIT_s0 .INIT=1'b1;
DFFC \u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_POWER_DOWN_s0  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n596_33 ),
	.CLK(I_sdrc_clk),
	.CLEAR(\u_sdrc_hs_top/n9_6 ),
	.Q(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_POWER_DOWN )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_POWER_DOWN_s0 .INIT=1'b0;
DFFC \u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_SELFREFRESH_s0  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n598_33 ),
	.CLK(I_sdrc_clk),
	.CLEAR(\u_sdrc_hs_top/n9_6 ),
	.Q(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_SELFREFRESH )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_SELFREFRESH_s0 .INIT=1'b0;
DFFC \u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_SELFREFRESH_WAIT_s0  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n602_32 ),
	.CLK(I_sdrc_clk),
	.CLEAR(\u_sdrc_hs_top/n9_6 ),
	.Q(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_SELFREFRESH_WAIT )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_SELFREFRESH_WAIT_s0 .INIT=1'b0;
DFFC \u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_SELFREFRESH_EXIT_s0  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n604_31 ),
	.CLK(I_sdrc_clk),
	.CLEAR(\u_sdrc_hs_top/n9_6 ),
	.Q(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_SELFREFRESH_EXIT )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_SELFREFRESH_EXIT_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_31_s0  (
	.D(IO_sdram_dq_in[31]),
	.CLK(I_sdrc_clk),
	.Q(O_sdrc_data[31])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_31_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_30_s0  (
	.D(IO_sdram_dq_in[30]),
	.CLK(I_sdrc_clk),
	.Q(O_sdrc_data[30])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_30_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_29_s0  (
	.D(IO_sdram_dq_in[29]),
	.CLK(I_sdrc_clk),
	.Q(O_sdrc_data[29])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_29_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_28_s0  (
	.D(IO_sdram_dq_in[28]),
	.CLK(I_sdrc_clk),
	.Q(O_sdrc_data[28])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_28_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_27_s0  (
	.D(IO_sdram_dq_in[27]),
	.CLK(I_sdrc_clk),
	.Q(O_sdrc_data[27])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_27_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_26_s0  (
	.D(IO_sdram_dq_in[26]),
	.CLK(I_sdrc_clk),
	.Q(O_sdrc_data[26])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_26_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_25_s0  (
	.D(IO_sdram_dq_in[25]),
	.CLK(I_sdrc_clk),
	.Q(O_sdrc_data[25])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_25_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_24_s0  (
	.D(IO_sdram_dq_in[24]),
	.CLK(I_sdrc_clk),
	.Q(O_sdrc_data[24])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_24_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_23_s0  (
	.D(IO_sdram_dq_in[23]),
	.CLK(I_sdrc_clk),
	.Q(O_sdrc_data[23])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_23_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_22_s0  (
	.D(IO_sdram_dq_in[22]),
	.CLK(I_sdrc_clk),
	.Q(O_sdrc_data[22])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_22_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_21_s0  (
	.D(IO_sdram_dq_in[21]),
	.CLK(I_sdrc_clk),
	.Q(O_sdrc_data[21])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_21_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_20_s0  (
	.D(IO_sdram_dq_in[20]),
	.CLK(I_sdrc_clk),
	.Q(O_sdrc_data[20])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_20_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_19_s0  (
	.D(IO_sdram_dq_in[19]),
	.CLK(I_sdrc_clk),
	.Q(O_sdrc_data[19])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_19_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_18_s0  (
	.D(IO_sdram_dq_in[18]),
	.CLK(I_sdrc_clk),
	.Q(O_sdrc_data[18])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_18_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_17_s0  (
	.D(IO_sdram_dq_in[17]),
	.CLK(I_sdrc_clk),
	.Q(O_sdrc_data[17])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_17_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_16_s0  (
	.D(IO_sdram_dq_in[16]),
	.CLK(I_sdrc_clk),
	.Q(O_sdrc_data[16])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_16_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_15_s0  (
	.D(IO_sdram_dq_in[15]),
	.CLK(I_sdrc_clk),
	.Q(O_sdrc_data[15])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_15_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_14_s0  (
	.D(IO_sdram_dq_in[14]),
	.CLK(I_sdrc_clk),
	.Q(O_sdrc_data[14])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_14_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_13_s0  (
	.D(IO_sdram_dq_in[13]),
	.CLK(I_sdrc_clk),
	.Q(O_sdrc_data[13])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_13_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_12_s0  (
	.D(IO_sdram_dq_in[12]),
	.CLK(I_sdrc_clk),
	.Q(O_sdrc_data[12])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_12_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_11_s0  (
	.D(IO_sdram_dq_in[11]),
	.CLK(I_sdrc_clk),
	.Q(O_sdrc_data[11])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_11_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_10_s0  (
	.D(IO_sdram_dq_in[10]),
	.CLK(I_sdrc_clk),
	.Q(O_sdrc_data[10])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_10_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_9_s0  (
	.D(IO_sdram_dq_in[9]),
	.CLK(I_sdrc_clk),
	.Q(O_sdrc_data[9])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_9_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_8_s0  (
	.D(IO_sdram_dq_in[8]),
	.CLK(I_sdrc_clk),
	.Q(O_sdrc_data[8])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_8_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_7_s0  (
	.D(IO_sdram_dq_in[7]),
	.CLK(I_sdrc_clk),
	.Q(O_sdrc_data[7])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_7_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_6_s0  (
	.D(IO_sdram_dq_in[6]),
	.CLK(I_sdrc_clk),
	.Q(O_sdrc_data[6])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_6_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_5_s0  (
	.D(IO_sdram_dq_in[5]),
	.CLK(I_sdrc_clk),
	.Q(O_sdrc_data[5])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_5_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_4_s0  (
	.D(IO_sdram_dq_in[4]),
	.CLK(I_sdrc_clk),
	.Q(O_sdrc_data[4])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_4_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_3_s0  (
	.D(IO_sdram_dq_in[3]),
	.CLK(I_sdrc_clk),
	.Q(O_sdrc_data[3])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_3_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_2_s0  (
	.D(IO_sdram_dq_in[2]),
	.CLK(I_sdrc_clk),
	.Q(O_sdrc_data[2])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_2_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_1_s0  (
	.D(IO_sdram_dq_in[1]),
	.CLK(I_sdrc_clk),
	.Q(O_sdrc_data[1])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_1_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_0_s0  (
	.D(IO_sdram_dq_in[0]),
	.CLK(I_sdrc_clk),
	.Q(O_sdrc_data[0])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_data_0_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_wen_n_s0  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n997_16 ),
	.CLK(I_sdrc_clk),
	.Q(\u_sdrc_hs_top/Sdram_wen_n )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_wen_n_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_cas_n_s0  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n1000_17 ),
	.CLK(I_sdrc_clk),
	.Q(\u_sdrc_hs_top/Sdram_cas_n )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_cas_n_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_ras_n_s0  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n1003_16 ),
	.CLK(I_sdrc_clk),
	.Q(\u_sdrc_hs_top/Sdram_ras_n )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_ras_n_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_ba_1_s0  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n1005_18 ),
	.CLK(I_sdrc_clk),
	.Q(\u_sdrc_hs_top/Sdram_ba [1])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_ba_1_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_ba_0_s0  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n1007_18 ),
	.CLK(I_sdrc_clk),
	.Q(\u_sdrc_hs_top/Sdram_ba [0])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_ba_0_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_addr_10_s0  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n1009_18 ),
	.CLK(I_sdrc_clk),
	.Q(\u_sdrc_hs_top/Sdram_addr [10])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_addr_10_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_addr_9_s0  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n1011_18 ),
	.CLK(I_sdrc_clk),
	.Q(\u_sdrc_hs_top/Sdram_addr [9])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_addr_9_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_addr_8_s0  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n1013_18 ),
	.CLK(I_sdrc_clk),
	.Q(\u_sdrc_hs_top/Sdram_addr [8])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_addr_8_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_addr_7_s0  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n1015_18 ),
	.CLK(I_sdrc_clk),
	.Q(\u_sdrc_hs_top/Sdram_addr [7])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_addr_7_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_addr_6_s0  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n1017_18 ),
	.CLK(I_sdrc_clk),
	.Q(\u_sdrc_hs_top/Sdram_addr [6])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_addr_6_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_addr_5_s0  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n1019_18 ),
	.CLK(I_sdrc_clk),
	.Q(\u_sdrc_hs_top/Sdram_addr [5])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_addr_5_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_addr_4_s0  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n1021_18 ),
	.CLK(I_sdrc_clk),
	.Q(\u_sdrc_hs_top/Sdram_addr [4])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_addr_4_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_addr_3_s0  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n1023_18 ),
	.CLK(I_sdrc_clk),
	.Q(\u_sdrc_hs_top/Sdram_addr [3])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_addr_3_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_addr_2_s0  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n1025_18 ),
	.CLK(I_sdrc_clk),
	.Q(\u_sdrc_hs_top/Sdram_addr [2])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_addr_2_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_addr_1_s0  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n1027_18 ),
	.CLK(I_sdrc_clk),
	.Q(\u_sdrc_hs_top/Sdram_addr [1])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_addr_1_s0 .INIT=1'b0;
DFF \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_addr_0_s0  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n1029_18 ),
	.CLK(I_sdrc_clk),
	.Q(\u_sdrc_hs_top/Sdram_addr [0])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_addr_0_s0 .INIT=1'b0;
DFFP \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_cs_n_s0  (
	.D(GND),
	.CLK(I_sdrc_clk),
	.PRESET(\u_sdrc_hs_top/n9_6 ),
	.Q(O_sdram_cs_n)
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_cs_n_s0 .INIT=1'b1;
DFFE \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd_7_s1  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n179_3 ),
	.CLK(I_sdrc_clk),
	.CE(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd_7_11 ),
	.Q(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd [7])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd_7_s1 .INIT=1'b0;
DFFE \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd_6_s1  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n180_3 ),
	.CLK(I_sdrc_clk),
	.CE(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd_7_11 ),
	.Q(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd [6])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd_6_s1 .INIT=1'b0;
DFFE \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd_5_s1  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n181_3 ),
	.CLK(I_sdrc_clk),
	.CE(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd_7_11 ),
	.Q(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd [5])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd_5_s1 .INIT=1'b0;
DFFE \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd_4_s1  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n182_3 ),
	.CLK(I_sdrc_clk),
	.CE(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd_7_11 ),
	.Q(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd [4])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd_4_s1 .INIT=1'b0;
DFFE \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd_3_s1  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n183_3 ),
	.CLK(I_sdrc_clk),
	.CE(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd_7_11 ),
	.Q(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd [3])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd_3_s1 .INIT=1'b0;
DFFE \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd_2_s1  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n184_3 ),
	.CLK(I_sdrc_clk),
	.CE(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd_7_11 ),
	.Q(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd [2])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd_2_s1 .INIT=1'b0;
DFFE \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd_1_s1  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n185_3 ),
	.CLK(I_sdrc_clk),
	.CE(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd_7_11 ),
	.Q(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd [1])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd_1_s1 .INIT=1'b0;
DFFE \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd_0_s1  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n186_3 ),
	.CLK(I_sdrc_clk),
	.CE(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd_7_11 ),
	.Q(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd [0])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_fsm_addr_col_wrd_0_s1 .INIT=1'b0;
(*gowin_io_reg = "FALSE" *) DFFCE \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_wr_data_valid_s1  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n759_8 ),
	.CLK(I_sdrc_clk),
	.CE(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_wr_data_valid_8 ),
	.CLEAR(\u_sdrc_hs_top/n9_6 ),
	.Q(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_wr_data_valid )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_wr_data_valid_s1 .INIT=1'b0;
DFFCE \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_cmd_ack_s4  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n80_31 ),
	.CLK(I_sdrc_clk),
	.CE(\u_sdrc_hs_top/u_sdrc_control_fsm/n80_29 ),
	.CLEAR(\u_sdrc_hs_top/n9_6 ),
	.Q(O_sdrc_cmd_ack)
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdrc_cmd_ack_s4 .INIT=1'b0;
DFFCE \u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num_8_s1  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n606_14 ),
	.CLK(I_sdrc_clk),
	.CE(\u_sdrc_hs_top/u_sdrc_control_fsm/n606_17 ),
	.CLEAR(\u_sdrc_hs_top/n9_6 ),
	.Q(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num [8])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num_8_s1 .INIT=1'b0;
DFFCE \u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num_7_s1  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n608_14 ),
	.CLK(I_sdrc_clk),
	.CE(\u_sdrc_hs_top/u_sdrc_control_fsm/n606_17 ),
	.CLEAR(\u_sdrc_hs_top/n9_6 ),
	.Q(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num [7])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num_7_s1 .INIT=1'b0;
DFFCE \u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num_6_s1  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n610_17 ),
	.CLK(I_sdrc_clk),
	.CE(\u_sdrc_hs_top/u_sdrc_control_fsm/n606_17 ),
	.CLEAR(\u_sdrc_hs_top/n9_6 ),
	.Q(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num [6])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num_6_s1 .INIT=1'b0;
DFFCE \u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num_5_s1  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n612_15 ),
	.CLK(I_sdrc_clk),
	.CE(\u_sdrc_hs_top/u_sdrc_control_fsm/n606_17 ),
	.CLEAR(\u_sdrc_hs_top/n9_6 ),
	.Q(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num [5])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num_5_s1 .INIT=1'b0;
DFFCE \u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num_4_s1  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n614_15 ),
	.CLK(I_sdrc_clk),
	.CE(\u_sdrc_hs_top/u_sdrc_control_fsm/n606_17 ),
	.CLEAR(\u_sdrc_hs_top/n9_6 ),
	.Q(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num [4])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num_4_s1 .INIT=1'b0;
DFFCE \u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num_3_s1  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n616_15 ),
	.CLK(I_sdrc_clk),
	.CE(\u_sdrc_hs_top/u_sdrc_control_fsm/n606_17 ),
	.CLEAR(\u_sdrc_hs_top/n9_6 ),
	.Q(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num [3])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num_3_s1 .INIT=1'b0;
DFFCE \u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num_2_s1  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n618_12 ),
	.CLK(I_sdrc_clk),
	.CE(\u_sdrc_hs_top/u_sdrc_control_fsm/n606_17 ),
	.CLEAR(\u_sdrc_hs_top/n9_6 ),
	.Q(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num [2])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num_2_s1 .INIT=1'b0;
DFFCE \u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num_1_s1  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n620_14 ),
	.CLK(I_sdrc_clk),
	.CE(\u_sdrc_hs_top/u_sdrc_control_fsm/n606_17 ),
	.CLEAR(\u_sdrc_hs_top/n9_6 ),
	.Q(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num [1])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num_1_s1 .INIT=1'b0;
DFFSE \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_cke_s3  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/Cmd_fsm_state.SDRC_STATE_DATAIN2ACTIVE ),
	.CLK(I_sdrc_clk),
	.CE(\u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_cke_7 ),
	.SET(\u_sdrc_hs_top/u_sdrc_control_fsm/n993_7 ),
	.Q(\u_sdrc_hs_top/Sdram_cke )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/O_sdram_cke_s3 .INIT=1'b1;
DFFC \u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num_0_s2  (
	.D(\u_sdrc_hs_top/u_sdrc_control_fsm/n622_17 ),
	.CLK(I_sdrc_clk),
	.CLEAR(\u_sdrc_hs_top/n9_6 ),
	.Q(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num [0])
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/Count_burst_num_0_s2 .INIT=1'b0;
INV \u_sdrc_hs_top/u_sdrc_control_fsm/IO_sdram_dq_0_s3  (
	.I(\u_sdrc_hs_top/u_sdrc_control_fsm/Ctrl_wr_data_valid ),
	.O(IO_sdram_dq_0_6)
);
LUT1 \u_sdrc_hs_top/u_sdrc_control_fsm/n87_s2  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay [0]),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n87_6 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n87_s2 .INIT=2'h1;
LUT1 \u_sdrc_hs_top/u_sdrc_control_fsm/n101_s2  (
	.I0(\u_sdrc_hs_top/u_sdrc_control_fsm/Count_cmd_delay2 [0]),
	.F(\u_sdrc_hs_top/u_sdrc_control_fsm/n101_6 )
);
defparam \u_sdrc_hs_top/u_sdrc_control_fsm/n101_s2 .INIT=2'h1;
endmodule
